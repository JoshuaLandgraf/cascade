// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

// Used with modifications by Joshua Landgraf

module cl_dma_pcis_slv
(
    input aclk,
    input aresetn,
    
    axi_bus_t.master sh_cl_dma_pcis_bus,
    axi_bus_t.master cl_axi_mstr_bus_1,
    axi_bus_t.master cl_axi_mstr_bus_2,
    axi_bus_t.master cl_axi_mstr_bus_3,
    axi_bus_t.master cl_axi_mstr_bus_4,
    
    axi_bus_t.slave lcl_cl_sh_ddra,
    axi_bus_t.slave lcl_cl_sh_ddrb,
    axi_bus_t.slave lcl_cl_sh_ddrd,
    
    axi_bus_t.slave cl_sh_ddr_bus
);

//----------------------------
// Internal signals
//----------------------------
axi_bus_t sh_cl_dma_pcis_q();
axi_bus_t cl_axi_mstr_bus_1_q();
axi_bus_t cl_axi_mstr_bus_2_q();
axi_bus_t cl_axi_mstr_bus_3_q();
axi_bus_t cl_axi_mstr_bus_4_q();
axi_bus_t cl_axi_mstr_bus_1_q2();
axi_bus_t cl_axi_mstr_bus_2_q2();
axi_bus_t cl_axi_mstr_bus_3_q2();
axi_bus_t cl_axi_mstr_bus_4_q2();
axi_bus_t cl_axi_mstr_bus_1_t();
axi_bus_t cl_axi_mstr_bus_2_t();
axi_bus_t cl_axi_mstr_bus_3_t();
axi_bus_t cl_axi_mstr_bus_4_t();
axi_bus_t lcl_cl_sh_ddra_q();
axi_bus_t lcl_cl_sh_ddrb_q();
axi_bus_t lcl_cl_sh_ddrd_q();
axi_bus_t lcl_cl_sh_ddra_q2();
axi_bus_t lcl_cl_sh_ddrb_q2();
axi_bus_t lcl_cl_sh_ddrd_q2();
axi_bus_t cl_sh_ddr_q();
axi_bus_t cl_sh_ddr_q2();
axi_bus_t sh_cl_pcis();

//----------------------------
// End Internal signals
//----------------------------


// Reset synchronizers
/*
(* dont_touch = "true" *) logic slr0_sync_aresetn;
(* dont_touch = "true" *) logic slr1_sync_aresetn;
(* dont_touch = "true" *) logic slr2_sync_aresetn;
lib_pipe #(.WIDTH(1), .STAGES(4)) SLR0_PIPE_RST_N (.clk(aclk), .rst_n(1'b1), .in_bus(aresetn), .out_bus(slr0_sync_aresetn));
lib_pipe #(.WIDTH(1), .STAGES(4)) SLR1_PIPE_RST_N (.clk(aclk), .rst_n(1'b1), .in_bus(aresetn), .out_bus(slr1_sync_aresetn));
lib_pipe #(.WIDTH(1), .STAGES(4)) SLR2_PIPE_RST_N (.clk(aclk), .rst_n(1'b1), .in_bus(aresetn), .out_bus(slr2_sync_aresetn));
*/

//----------------------------
// flop the dma_pcis interface input of CL
//----------------------------

// AXI4 Register Slice for dma_pcis interface
axi_register_slice PCI_AXL_REG_SLC_1 (
    .aclk          (aclk),
    .aresetn       (aresetn),
    .s_axi_awid    (sh_cl_dma_pcis_bus.awid),
    .s_axi_awaddr  (sh_cl_dma_pcis_bus.awaddr),
    .s_axi_awlen   (sh_cl_dma_pcis_bus.awlen),
    .s_axi_awvalid (sh_cl_dma_pcis_bus.awvalid),
    .s_axi_awsize  (sh_cl_dma_pcis_bus.awsize),
    .s_axi_awready (sh_cl_dma_pcis_bus.awready),
    .s_axi_wdata   (sh_cl_dma_pcis_bus.wdata),
    .s_axi_wstrb   (sh_cl_dma_pcis_bus.wstrb),
    .s_axi_wlast   (sh_cl_dma_pcis_bus.wlast),
    .s_axi_wvalid  (sh_cl_dma_pcis_bus.wvalid),
    .s_axi_wready  (sh_cl_dma_pcis_bus.wready),
    .s_axi_bid     (sh_cl_dma_pcis_bus.bid),
    .s_axi_bresp   (sh_cl_dma_pcis_bus.bresp),
    .s_axi_bvalid  (sh_cl_dma_pcis_bus.bvalid),
    .s_axi_bready  (sh_cl_dma_pcis_bus.bready),
    .s_axi_arid    (sh_cl_dma_pcis_bus.arid),
    .s_axi_araddr  (sh_cl_dma_pcis_bus.araddr),
    .s_axi_arlen   (sh_cl_dma_pcis_bus.arlen),
    .s_axi_arvalid (sh_cl_dma_pcis_bus.arvalid),
    .s_axi_arsize  (sh_cl_dma_pcis_bus.arsize),
    .s_axi_arready (sh_cl_dma_pcis_bus.arready),
    .s_axi_rid     (sh_cl_dma_pcis_bus.rid),
    .s_axi_rdata   (sh_cl_dma_pcis_bus.rdata),
    .s_axi_rresp   (sh_cl_dma_pcis_bus.rresp),
    .s_axi_rlast   (sh_cl_dma_pcis_bus.rlast),
    .s_axi_rvalid  (sh_cl_dma_pcis_bus.rvalid),
    .s_axi_rready  (sh_cl_dma_pcis_bus.rready),
    
    .m_axi_awid    (sh_cl_dma_pcis_q.awid),
    .m_axi_awaddr  (sh_cl_dma_pcis_q.awaddr),
    .m_axi_awlen   (sh_cl_dma_pcis_q.awlen),
    .m_axi_awvalid (sh_cl_dma_pcis_q.awvalid),
    .m_axi_awsize  (sh_cl_dma_pcis_q.awsize),
    .m_axi_awready (sh_cl_dma_pcis_q.awready),
    .m_axi_wdata   (sh_cl_dma_pcis_q.wdata),
    .m_axi_wstrb   (sh_cl_dma_pcis_q.wstrb),
    .m_axi_wvalid  (sh_cl_dma_pcis_q.wvalid),
    .m_axi_wlast   (sh_cl_dma_pcis_q.wlast),
    .m_axi_wready  (sh_cl_dma_pcis_q.wready),
    .m_axi_bresp   (sh_cl_dma_pcis_q.bresp),
    .m_axi_bvalid  (sh_cl_dma_pcis_q.bvalid),
    .m_axi_bid     (sh_cl_dma_pcis_q.bid),
    .m_axi_bready  (sh_cl_dma_pcis_q.bready),
    .m_axi_arid    (sh_cl_dma_pcis_q.arid),
    .m_axi_araddr  (sh_cl_dma_pcis_q.araddr),
    .m_axi_arlen   (sh_cl_dma_pcis_q.arlen),
    .m_axi_arsize  (sh_cl_dma_pcis_q.arsize),
    .m_axi_arvalid (sh_cl_dma_pcis_q.arvalid),
    .m_axi_arready (sh_cl_dma_pcis_q.arready),
    .m_axi_rid     (sh_cl_dma_pcis_q.rid),
    .m_axi_rdata   (sh_cl_dma_pcis_q.rdata),
    .m_axi_rresp   (sh_cl_dma_pcis_q.rresp),
    .m_axi_rlast   (sh_cl_dma_pcis_q.rlast),
    .m_axi_rvalid  (sh_cl_dma_pcis_q.rvalid),
    .m_axi_rready  (sh_cl_dma_pcis_q.rready)
);

//-----------------------------------------------------
// tie-off unused signals to prevent critical warnings
//-----------------------------------------------------
assign sh_cl_dma_pcis_q.rid[15:6] = 10'b0;
assign sh_cl_dma_pcis_q.bid[15:6] = 10'b0;

//----------------------------
// flop the master interfaces input of CL
//----------------------------
axi_register_slice MSTR_1_AXL_REG_SLC_1 (
    .aclk          (aclk),
    .aresetn       (aresetn),
    .s_axi_awid    (cl_axi_mstr_bus_1.awid),
    .s_axi_awaddr  (cl_axi_mstr_bus_1.awaddr),
    .s_axi_awlen   (cl_axi_mstr_bus_1.awlen),
    .s_axi_awvalid (cl_axi_mstr_bus_1.awvalid),
    .s_axi_awsize  (cl_axi_mstr_bus_1.awsize),
    .s_axi_awready (cl_axi_mstr_bus_1.awready),
    .s_axi_wdata   (cl_axi_mstr_bus_1.wdata),
    .s_axi_wstrb   (cl_axi_mstr_bus_1.wstrb),
    .s_axi_wlast   (cl_axi_mstr_bus_1.wlast),
    .s_axi_wvalid  (cl_axi_mstr_bus_1.wvalid),
    .s_axi_wready  (cl_axi_mstr_bus_1.wready),
    .s_axi_bid     (cl_axi_mstr_bus_1.bid),
    .s_axi_bresp   (cl_axi_mstr_bus_1.bresp),
    .s_axi_bvalid  (cl_axi_mstr_bus_1.bvalid),
    .s_axi_bready  (cl_axi_mstr_bus_1.bready),
    .s_axi_arid    (cl_axi_mstr_bus_1.arid),
    .s_axi_araddr  (cl_axi_mstr_bus_1.araddr),
    .s_axi_arlen   (cl_axi_mstr_bus_1.arlen),
    .s_axi_arvalid (cl_axi_mstr_bus_1.arvalid),
    .s_axi_arsize  (cl_axi_mstr_bus_1.arsize),
    .s_axi_arready (cl_axi_mstr_bus_1.arready),
    .s_axi_rid     (cl_axi_mstr_bus_1.rid),
    .s_axi_rdata   (cl_axi_mstr_bus_1.rdata),
    .s_axi_rresp   (cl_axi_mstr_bus_1.rresp),
    .s_axi_rlast   (cl_axi_mstr_bus_1.rlast),
    .s_axi_rvalid  (cl_axi_mstr_bus_1.rvalid),
    .s_axi_rready  (cl_axi_mstr_bus_1.rready),
    
    .m_axi_awid    (cl_axi_mstr_bus_1_q.awid),
    .m_axi_awaddr  (cl_axi_mstr_bus_1_q.awaddr),
    .m_axi_awlen   (cl_axi_mstr_bus_1_q.awlen),
    .m_axi_awvalid (cl_axi_mstr_bus_1_q.awvalid),
    .m_axi_awsize  (cl_axi_mstr_bus_1_q.awsize),
    .m_axi_awready (cl_axi_mstr_bus_1_q.awready),
    .m_axi_wdata   (cl_axi_mstr_bus_1_q.wdata),
    .m_axi_wstrb   (cl_axi_mstr_bus_1_q.wstrb),
    .m_axi_wvalid  (cl_axi_mstr_bus_1_q.wvalid),
    .m_axi_wlast   (cl_axi_mstr_bus_1_q.wlast),
    .m_axi_wready  (cl_axi_mstr_bus_1_q.wready),
    .m_axi_bresp   (cl_axi_mstr_bus_1_q.bresp),
    .m_axi_bvalid  (cl_axi_mstr_bus_1_q.bvalid),
    .m_axi_bid     (cl_axi_mstr_bus_1_q.bid),
    .m_axi_bready  (cl_axi_mstr_bus_1_q.bready),
    .m_axi_arid    (cl_axi_mstr_bus_1_q.arid),
    .m_axi_araddr  (cl_axi_mstr_bus_1_q.araddr),
    .m_axi_arlen   (cl_axi_mstr_bus_1_q.arlen),
    .m_axi_arsize  (cl_axi_mstr_bus_1_q.arsize),
    .m_axi_arvalid (cl_axi_mstr_bus_1_q.arvalid),
    .m_axi_arready (cl_axi_mstr_bus_1_q.arready),
    .m_axi_rid     (cl_axi_mstr_bus_1_q.rid),
    .m_axi_rdata   (cl_axi_mstr_bus_1_q.rdata),
    .m_axi_rresp   (cl_axi_mstr_bus_1_q.rresp),
    .m_axi_rlast   (cl_axi_mstr_bus_1_q.rlast),
    .m_axi_rvalid  (cl_axi_mstr_bus_1_q.rvalid),
    .m_axi_rready  (cl_axi_mstr_bus_1_q.rready)
);
axi_register_slice MSTR_1_AXL_REG_SLC_2 (
    .aclk          (aclk),
    .aresetn       (aresetn),
    .s_axi_awid    (cl_axi_mstr_bus_1_q.awid),
    .s_axi_awaddr  (cl_axi_mstr_bus_1_q.awaddr),
    .s_axi_awlen   (cl_axi_mstr_bus_1_q.awlen),
    .s_axi_awvalid (cl_axi_mstr_bus_1_q.awvalid),
    .s_axi_awsize  (cl_axi_mstr_bus_1_q.awsize),
    .s_axi_awready (cl_axi_mstr_bus_1_q.awready),
    .s_axi_wdata   (cl_axi_mstr_bus_1_q.wdata),
    .s_axi_wstrb   (cl_axi_mstr_bus_1_q.wstrb),
    .s_axi_wlast   (cl_axi_mstr_bus_1_q.wlast),
    .s_axi_wvalid  (cl_axi_mstr_bus_1_q.wvalid),
    .s_axi_wready  (cl_axi_mstr_bus_1_q.wready),
    .s_axi_bid     (cl_axi_mstr_bus_1_q.bid),
    .s_axi_bresp   (cl_axi_mstr_bus_1_q.bresp),
    .s_axi_bvalid  (cl_axi_mstr_bus_1_q.bvalid),
    .s_axi_bready  (cl_axi_mstr_bus_1_q.bready),
    .s_axi_arid    (cl_axi_mstr_bus_1_q.arid),
    .s_axi_araddr  (cl_axi_mstr_bus_1_q.araddr),
    .s_axi_arlen   (cl_axi_mstr_bus_1_q.arlen),
    .s_axi_arvalid (cl_axi_mstr_bus_1_q.arvalid),
    .s_axi_arsize  (cl_axi_mstr_bus_1_q.arsize),
    .s_axi_arready (cl_axi_mstr_bus_1_q.arready),
    .s_axi_rid     (cl_axi_mstr_bus_1_q.rid),
    .s_axi_rdata   (cl_axi_mstr_bus_1_q.rdata),
    .s_axi_rresp   (cl_axi_mstr_bus_1_q.rresp),
    .s_axi_rlast   (cl_axi_mstr_bus_1_q.rlast),
    .s_axi_rvalid  (cl_axi_mstr_bus_1_q.rvalid),
    .s_axi_rready  (cl_axi_mstr_bus_1_q.rready),
    
    .m_axi_awid    (cl_axi_mstr_bus_1_q2.awid),
    .m_axi_awaddr  (cl_axi_mstr_bus_1_q2.awaddr),
    .m_axi_awlen   (cl_axi_mstr_bus_1_q2.awlen),
    .m_axi_awvalid (cl_axi_mstr_bus_1_q2.awvalid),
    .m_axi_awsize  (cl_axi_mstr_bus_1_q2.awsize),
    .m_axi_awready (cl_axi_mstr_bus_1_q2.awready),
    .m_axi_wdata   (cl_axi_mstr_bus_1_q2.wdata),
    .m_axi_wstrb   (cl_axi_mstr_bus_1_q2.wstrb),
    .m_axi_wvalid  (cl_axi_mstr_bus_1_q2.wvalid),
    .m_axi_wlast   (cl_axi_mstr_bus_1_q2.wlast),
    .m_axi_wready  (cl_axi_mstr_bus_1_q2.wready),
    .m_axi_bresp   (cl_axi_mstr_bus_1_q2.bresp),
    .m_axi_bvalid  (cl_axi_mstr_bus_1_q2.bvalid),
    .m_axi_bid     (cl_axi_mstr_bus_1_q2.bid),
    .m_axi_bready  (cl_axi_mstr_bus_1_q2.bready),
    .m_axi_arid    (cl_axi_mstr_bus_1_q2.arid),
    .m_axi_araddr  (cl_axi_mstr_bus_1_q2.araddr),
    .m_axi_arlen   (cl_axi_mstr_bus_1_q2.arlen),
    .m_axi_arsize  (cl_axi_mstr_bus_1_q2.arsize),
    .m_axi_arvalid (cl_axi_mstr_bus_1_q2.arvalid),
    .m_axi_arready (cl_axi_mstr_bus_1_q2.arready),
    .m_axi_rid     (cl_axi_mstr_bus_1_q2.rid),
    .m_axi_rdata   (cl_axi_mstr_bus_1_q2.rdata),
    .m_axi_rresp   (cl_axi_mstr_bus_1_q2.rresp),
    .m_axi_rlast   (cl_axi_mstr_bus_1_q2.rlast),
    .m_axi_rvalid  (cl_axi_mstr_bus_1_q2.rvalid),
    .m_axi_rready  (cl_axi_mstr_bus_1_q2.rready)
);
axi_register_slice MSTR_2_AXL_REG_SLC_1 (
    .aclk          (aclk),
    .aresetn       (aresetn),
    .s_axi_awid    (cl_axi_mstr_bus_2.awid),
    .s_axi_awaddr  (cl_axi_mstr_bus_2.awaddr),
    .s_axi_awlen   (cl_axi_mstr_bus_2.awlen),
    .s_axi_awvalid (cl_axi_mstr_bus_2.awvalid),
    .s_axi_awsize  (cl_axi_mstr_bus_2.awsize),
    .s_axi_awready (cl_axi_mstr_bus_2.awready),
    .s_axi_wdata   (cl_axi_mstr_bus_2.wdata),
    .s_axi_wstrb   (cl_axi_mstr_bus_2.wstrb),
    .s_axi_wlast   (cl_axi_mstr_bus_2.wlast),
    .s_axi_wvalid  (cl_axi_mstr_bus_2.wvalid),
    .s_axi_wready  (cl_axi_mstr_bus_2.wready),
    .s_axi_bid     (cl_axi_mstr_bus_2.bid),
    .s_axi_bresp   (cl_axi_mstr_bus_2.bresp),
    .s_axi_bvalid  (cl_axi_mstr_bus_2.bvalid),
    .s_axi_bready  (cl_axi_mstr_bus_2.bready),
    .s_axi_arid    (cl_axi_mstr_bus_2.arid),
    .s_axi_araddr  (cl_axi_mstr_bus_2.araddr),
    .s_axi_arlen   (cl_axi_mstr_bus_2.arlen),
    .s_axi_arvalid (cl_axi_mstr_bus_2.arvalid),
    .s_axi_arsize  (cl_axi_mstr_bus_2.arsize),
    .s_axi_arready (cl_axi_mstr_bus_2.arready),
    .s_axi_rid     (cl_axi_mstr_bus_2.rid),
    .s_axi_rdata   (cl_axi_mstr_bus_2.rdata),
    .s_axi_rresp   (cl_axi_mstr_bus_2.rresp),
    .s_axi_rlast   (cl_axi_mstr_bus_2.rlast),
    .s_axi_rvalid  (cl_axi_mstr_bus_2.rvalid),
    .s_axi_rready  (cl_axi_mstr_bus_2.rready),
    
    .m_axi_awid    (cl_axi_mstr_bus_2_q.awid),
    .m_axi_awaddr  (cl_axi_mstr_bus_2_q.awaddr),
    .m_axi_awlen   (cl_axi_mstr_bus_2_q.awlen),
    .m_axi_awvalid (cl_axi_mstr_bus_2_q.awvalid),
    .m_axi_awsize  (cl_axi_mstr_bus_2_q.awsize),
    .m_axi_awready (cl_axi_mstr_bus_2_q.awready),
    .m_axi_wdata   (cl_axi_mstr_bus_2_q.wdata),
    .m_axi_wstrb   (cl_axi_mstr_bus_2_q.wstrb),
    .m_axi_wvalid  (cl_axi_mstr_bus_2_q.wvalid),
    .m_axi_wlast   (cl_axi_mstr_bus_2_q.wlast),
    .m_axi_wready  (cl_axi_mstr_bus_2_q.wready),
    .m_axi_bresp   (cl_axi_mstr_bus_2_q.bresp),
    .m_axi_bvalid  (cl_axi_mstr_bus_2_q.bvalid),
    .m_axi_bid     (cl_axi_mstr_bus_2_q.bid),
    .m_axi_bready  (cl_axi_mstr_bus_2_q.bready),
    .m_axi_arid    (cl_axi_mstr_bus_2_q.arid),
    .m_axi_araddr  (cl_axi_mstr_bus_2_q.araddr),
    .m_axi_arlen   (cl_axi_mstr_bus_2_q.arlen),
    .m_axi_arsize  (cl_axi_mstr_bus_2_q.arsize),
    .m_axi_arvalid (cl_axi_mstr_bus_2_q.arvalid),
    .m_axi_arready (cl_axi_mstr_bus_2_q.arready),
    .m_axi_rid     (cl_axi_mstr_bus_2_q.rid),
    .m_axi_rdata   (cl_axi_mstr_bus_2_q.rdata),
    .m_axi_rresp   (cl_axi_mstr_bus_2_q.rresp),
    .m_axi_rlast   (cl_axi_mstr_bus_2_q.rlast),
    .m_axi_rvalid  (cl_axi_mstr_bus_2_q.rvalid),
    .m_axi_rready  (cl_axi_mstr_bus_2_q.rready)
);
axi_register_slice MSTR_2_AXL_REG_SLC_2 (
    .aclk          (aclk),
    .aresetn       (aresetn),
    .s_axi_awid    (cl_axi_mstr_bus_2_q.awid),
    .s_axi_awaddr  (cl_axi_mstr_bus_2_q.awaddr),
    .s_axi_awlen   (cl_axi_mstr_bus_2_q.awlen),
    .s_axi_awvalid (cl_axi_mstr_bus_2_q.awvalid),
    .s_axi_awsize  (cl_axi_mstr_bus_2_q.awsize),
    .s_axi_awready (cl_axi_mstr_bus_2_q.awready),
    .s_axi_wdata   (cl_axi_mstr_bus_2_q.wdata),
    .s_axi_wstrb   (cl_axi_mstr_bus_2_q.wstrb),
    .s_axi_wlast   (cl_axi_mstr_bus_2_q.wlast),
    .s_axi_wvalid  (cl_axi_mstr_bus_2_q.wvalid),
    .s_axi_wready  (cl_axi_mstr_bus_2_q.wready),
    .s_axi_bid     (cl_axi_mstr_bus_2_q.bid),
    .s_axi_bresp   (cl_axi_mstr_bus_2_q.bresp),
    .s_axi_bvalid  (cl_axi_mstr_bus_2_q.bvalid),
    .s_axi_bready  (cl_axi_mstr_bus_2_q.bready),
    .s_axi_arid    (cl_axi_mstr_bus_2_q.arid),
    .s_axi_araddr  (cl_axi_mstr_bus_2_q.araddr),
    .s_axi_arlen   (cl_axi_mstr_bus_2_q.arlen),
    .s_axi_arvalid (cl_axi_mstr_bus_2_q.arvalid),
    .s_axi_arsize  (cl_axi_mstr_bus_2_q.arsize),
    .s_axi_arready (cl_axi_mstr_bus_2_q.arready),
    .s_axi_rid     (cl_axi_mstr_bus_2_q.rid),
    .s_axi_rdata   (cl_axi_mstr_bus_2_q.rdata),
    .s_axi_rresp   (cl_axi_mstr_bus_2_q.rresp),
    .s_axi_rlast   (cl_axi_mstr_bus_2_q.rlast),
    .s_axi_rvalid  (cl_axi_mstr_bus_2_q.rvalid),
    .s_axi_rready  (cl_axi_mstr_bus_2_q.rready),
    
    .m_axi_awid    (cl_axi_mstr_bus_2_q2.awid),
    .m_axi_awaddr  (cl_axi_mstr_bus_2_q2.awaddr),
    .m_axi_awlen   (cl_axi_mstr_bus_2_q2.awlen),
    .m_axi_awvalid (cl_axi_mstr_bus_2_q2.awvalid),
    .m_axi_awsize  (cl_axi_mstr_bus_2_q2.awsize),
    .m_axi_awready (cl_axi_mstr_bus_2_q2.awready),
    .m_axi_wdata   (cl_axi_mstr_bus_2_q2.wdata),
    .m_axi_wstrb   (cl_axi_mstr_bus_2_q2.wstrb),
    .m_axi_wvalid  (cl_axi_mstr_bus_2_q2.wvalid),
    .m_axi_wlast   (cl_axi_mstr_bus_2_q2.wlast),
    .m_axi_wready  (cl_axi_mstr_bus_2_q2.wready),
    .m_axi_bresp   (cl_axi_mstr_bus_2_q2.bresp),
    .m_axi_bvalid  (cl_axi_mstr_bus_2_q2.bvalid),
    .m_axi_bid     (cl_axi_mstr_bus_2_q2.bid),
    .m_axi_bready  (cl_axi_mstr_bus_2_q2.bready),
    .m_axi_arid    (cl_axi_mstr_bus_2_q2.arid),
    .m_axi_araddr  (cl_axi_mstr_bus_2_q2.araddr),
    .m_axi_arlen   (cl_axi_mstr_bus_2_q2.arlen),
    .m_axi_arsize  (cl_axi_mstr_bus_2_q2.arsize),
    .m_axi_arvalid (cl_axi_mstr_bus_2_q2.arvalid),
    .m_axi_arready (cl_axi_mstr_bus_2_q2.arready),
    .m_axi_rid     (cl_axi_mstr_bus_2_q2.rid),
    .m_axi_rdata   (cl_axi_mstr_bus_2_q2.rdata),
    .m_axi_rresp   (cl_axi_mstr_bus_2_q2.rresp),
    .m_axi_rlast   (cl_axi_mstr_bus_2_q2.rlast),
    .m_axi_rvalid  (cl_axi_mstr_bus_2_q2.rvalid),
    .m_axi_rready  (cl_axi_mstr_bus_2_q2.rready)
);
axi_register_slice MSTR_3_AXL_REG_SLC_1 (
    .aclk          (aclk),
    .aresetn       (aresetn),
    .s_axi_awid    (cl_axi_mstr_bus_3.awid),
    .s_axi_awaddr  (cl_axi_mstr_bus_3.awaddr),
    .s_axi_awlen   (cl_axi_mstr_bus_3.awlen),
    .s_axi_awvalid (cl_axi_mstr_bus_3.awvalid),
    .s_axi_awsize  (cl_axi_mstr_bus_3.awsize),
    .s_axi_awready (cl_axi_mstr_bus_3.awready),
    .s_axi_wdata   (cl_axi_mstr_bus_3.wdata),
    .s_axi_wstrb   (cl_axi_mstr_bus_3.wstrb),
    .s_axi_wlast   (cl_axi_mstr_bus_3.wlast),
    .s_axi_wvalid  (cl_axi_mstr_bus_3.wvalid),
    .s_axi_wready  (cl_axi_mstr_bus_3.wready),
    .s_axi_bid     (cl_axi_mstr_bus_3.bid),
    .s_axi_bresp   (cl_axi_mstr_bus_3.bresp),
    .s_axi_bvalid  (cl_axi_mstr_bus_3.bvalid),
    .s_axi_bready  (cl_axi_mstr_bus_3.bready),
    .s_axi_arid    (cl_axi_mstr_bus_3.arid),
    .s_axi_araddr  (cl_axi_mstr_bus_3.araddr),
    .s_axi_arlen   (cl_axi_mstr_bus_3.arlen),
    .s_axi_arvalid (cl_axi_mstr_bus_3.arvalid),
    .s_axi_arsize  (cl_axi_mstr_bus_3.arsize),
    .s_axi_arready (cl_axi_mstr_bus_3.arready),
    .s_axi_rid     (cl_axi_mstr_bus_3.rid),
    .s_axi_rdata   (cl_axi_mstr_bus_3.rdata),
    .s_axi_rresp   (cl_axi_mstr_bus_3.rresp),
    .s_axi_rlast   (cl_axi_mstr_bus_3.rlast),
    .s_axi_rvalid  (cl_axi_mstr_bus_3.rvalid),
    .s_axi_rready  (cl_axi_mstr_bus_3.rready),
    
    .m_axi_awid    (cl_axi_mstr_bus_3_q.awid),
    .m_axi_awaddr  (cl_axi_mstr_bus_3_q.awaddr),
    .m_axi_awlen   (cl_axi_mstr_bus_3_q.awlen),
    .m_axi_awvalid (cl_axi_mstr_bus_3_q.awvalid),
    .m_axi_awsize  (cl_axi_mstr_bus_3_q.awsize),
    .m_axi_awready (cl_axi_mstr_bus_3_q.awready),
    .m_axi_wdata   (cl_axi_mstr_bus_3_q.wdata),
    .m_axi_wstrb   (cl_axi_mstr_bus_3_q.wstrb),
    .m_axi_wvalid  (cl_axi_mstr_bus_3_q.wvalid),
    .m_axi_wlast   (cl_axi_mstr_bus_3_q.wlast),
    .m_axi_wready  (cl_axi_mstr_bus_3_q.wready),
    .m_axi_bresp   (cl_axi_mstr_bus_3_q.bresp),
    .m_axi_bvalid  (cl_axi_mstr_bus_3_q.bvalid),
    .m_axi_bid     (cl_axi_mstr_bus_3_q.bid),
    .m_axi_bready  (cl_axi_mstr_bus_3_q.bready),
    .m_axi_arid    (cl_axi_mstr_bus_3_q.arid),
    .m_axi_araddr  (cl_axi_mstr_bus_3_q.araddr),
    .m_axi_arlen   (cl_axi_mstr_bus_3_q.arlen),
    .m_axi_arsize  (cl_axi_mstr_bus_3_q.arsize),
    .m_axi_arvalid (cl_axi_mstr_bus_3_q.arvalid),
    .m_axi_arready (cl_axi_mstr_bus_3_q.arready),
    .m_axi_rid     (cl_axi_mstr_bus_3_q.rid),
    .m_axi_rdata   (cl_axi_mstr_bus_3_q.rdata),
    .m_axi_rresp   (cl_axi_mstr_bus_3_q.rresp),
    .m_axi_rlast   (cl_axi_mstr_bus_3_q.rlast),
    .m_axi_rvalid  (cl_axi_mstr_bus_3_q.rvalid),
    .m_axi_rready  (cl_axi_mstr_bus_3_q.rready)
);
axi_register_slice MSTR_3_AXL_REG_SLC_2 (
    .aclk          (aclk),
    .aresetn       (aresetn),
    .s_axi_awid    (cl_axi_mstr_bus_3_q.awid),
    .s_axi_awaddr  (cl_axi_mstr_bus_3_q.awaddr),
    .s_axi_awlen   (cl_axi_mstr_bus_3_q.awlen),
    .s_axi_awvalid (cl_axi_mstr_bus_3_q.awvalid),
    .s_axi_awsize  (cl_axi_mstr_bus_3_q.awsize),
    .s_axi_awready (cl_axi_mstr_bus_3_q.awready),
    .s_axi_wdata   (cl_axi_mstr_bus_3_q.wdata),
    .s_axi_wstrb   (cl_axi_mstr_bus_3_q.wstrb),
    .s_axi_wlast   (cl_axi_mstr_bus_3_q.wlast),
    .s_axi_wvalid  (cl_axi_mstr_bus_3_q.wvalid),
    .s_axi_wready  (cl_axi_mstr_bus_3_q.wready),
    .s_axi_bid     (cl_axi_mstr_bus_3_q.bid),
    .s_axi_bresp   (cl_axi_mstr_bus_3_q.bresp),
    .s_axi_bvalid  (cl_axi_mstr_bus_3_q.bvalid),
    .s_axi_bready  (cl_axi_mstr_bus_3_q.bready),
    .s_axi_arid    (cl_axi_mstr_bus_3_q.arid),
    .s_axi_araddr  (cl_axi_mstr_bus_3_q.araddr),
    .s_axi_arlen   (cl_axi_mstr_bus_3_q.arlen),
    .s_axi_arvalid (cl_axi_mstr_bus_3_q.arvalid),
    .s_axi_arsize  (cl_axi_mstr_bus_3_q.arsize),
    .s_axi_arready (cl_axi_mstr_bus_3_q.arready),
    .s_axi_rid     (cl_axi_mstr_bus_3_q.rid),
    .s_axi_rdata   (cl_axi_mstr_bus_3_q.rdata),
    .s_axi_rresp   (cl_axi_mstr_bus_3_q.rresp),
    .s_axi_rlast   (cl_axi_mstr_bus_3_q.rlast),
    .s_axi_rvalid  (cl_axi_mstr_bus_3_q.rvalid),
    .s_axi_rready  (cl_axi_mstr_bus_3_q.rready),
    
    .m_axi_awid    (cl_axi_mstr_bus_3_q2.awid),
    .m_axi_awaddr  (cl_axi_mstr_bus_3_q2.awaddr),
    .m_axi_awlen   (cl_axi_mstr_bus_3_q2.awlen),
    .m_axi_awvalid (cl_axi_mstr_bus_3_q2.awvalid),
    .m_axi_awsize  (cl_axi_mstr_bus_3_q2.awsize),
    .m_axi_awready (cl_axi_mstr_bus_3_q2.awready),
    .m_axi_wdata   (cl_axi_mstr_bus_3_q2.wdata),
    .m_axi_wstrb   (cl_axi_mstr_bus_3_q2.wstrb),
    .m_axi_wvalid  (cl_axi_mstr_bus_3_q2.wvalid),
    .m_axi_wlast   (cl_axi_mstr_bus_3_q2.wlast),
    .m_axi_wready  (cl_axi_mstr_bus_3_q2.wready),
    .m_axi_bresp   (cl_axi_mstr_bus_3_q2.bresp),
    .m_axi_bvalid  (cl_axi_mstr_bus_3_q2.bvalid),
    .m_axi_bid     (cl_axi_mstr_bus_3_q2.bid),
    .m_axi_bready  (cl_axi_mstr_bus_3_q2.bready),
    .m_axi_arid    (cl_axi_mstr_bus_3_q2.arid),
    .m_axi_araddr  (cl_axi_mstr_bus_3_q2.araddr),
    .m_axi_arlen   (cl_axi_mstr_bus_3_q2.arlen),
    .m_axi_arsize  (cl_axi_mstr_bus_3_q2.arsize),
    .m_axi_arvalid (cl_axi_mstr_bus_3_q2.arvalid),
    .m_axi_arready (cl_axi_mstr_bus_3_q2.arready),
    .m_axi_rid     (cl_axi_mstr_bus_3_q2.rid),
    .m_axi_rdata   (cl_axi_mstr_bus_3_q2.rdata),
    .m_axi_rresp   (cl_axi_mstr_bus_3_q2.rresp),
    .m_axi_rlast   (cl_axi_mstr_bus_3_q2.rlast),
    .m_axi_rvalid  (cl_axi_mstr_bus_3_q2.rvalid),
    .m_axi_rready  (cl_axi_mstr_bus_3_q2.rready)
);
axi_register_slice MSTR_4_AXL_REG_SLC_1 (
    .aclk          (aclk),
    .aresetn       (aresetn),
    .s_axi_awid    (cl_axi_mstr_bus_4.awid),
    .s_axi_awaddr  (cl_axi_mstr_bus_4.awaddr),
    .s_axi_awlen   (cl_axi_mstr_bus_4.awlen),
    .s_axi_awvalid (cl_axi_mstr_bus_4.awvalid),
    .s_axi_awsize  (cl_axi_mstr_bus_4.awsize),
    .s_axi_awready (cl_axi_mstr_bus_4.awready),
    .s_axi_wdata   (cl_axi_mstr_bus_4.wdata),
    .s_axi_wstrb   (cl_axi_mstr_bus_4.wstrb),
    .s_axi_wlast   (cl_axi_mstr_bus_4.wlast),
    .s_axi_wvalid  (cl_axi_mstr_bus_4.wvalid),
    .s_axi_wready  (cl_axi_mstr_bus_4.wready),
    .s_axi_bid     (cl_axi_mstr_bus_4.bid),
    .s_axi_bresp   (cl_axi_mstr_bus_4.bresp),
    .s_axi_bvalid  (cl_axi_mstr_bus_4.bvalid),
    .s_axi_bready  (cl_axi_mstr_bus_4.bready),
    .s_axi_arid    (cl_axi_mstr_bus_4.arid),
    .s_axi_araddr  (cl_axi_mstr_bus_4.araddr),
    .s_axi_arlen   (cl_axi_mstr_bus_4.arlen),
    .s_axi_arvalid (cl_axi_mstr_bus_4.arvalid),
    .s_axi_arsize  (cl_axi_mstr_bus_4.arsize),
    .s_axi_arready (cl_axi_mstr_bus_4.arready),
    .s_axi_rid     (cl_axi_mstr_bus_4.rid),
    .s_axi_rdata   (cl_axi_mstr_bus_4.rdata),
    .s_axi_rresp   (cl_axi_mstr_bus_4.rresp),
    .s_axi_rlast   (cl_axi_mstr_bus_4.rlast),
    .s_axi_rvalid  (cl_axi_mstr_bus_4.rvalid),
    .s_axi_rready  (cl_axi_mstr_bus_4.rready),
    
    .m_axi_awid    (cl_axi_mstr_bus_4_q.awid),
    .m_axi_awaddr  (cl_axi_mstr_bus_4_q.awaddr),
    .m_axi_awlen   (cl_axi_mstr_bus_4_q.awlen),
    .m_axi_awvalid (cl_axi_mstr_bus_4_q.awvalid),
    .m_axi_awsize  (cl_axi_mstr_bus_4_q.awsize),
    .m_axi_awready (cl_axi_mstr_bus_4_q.awready),
    .m_axi_wdata   (cl_axi_mstr_bus_4_q.wdata),
    .m_axi_wstrb   (cl_axi_mstr_bus_4_q.wstrb),
    .m_axi_wvalid  (cl_axi_mstr_bus_4_q.wvalid),
    .m_axi_wlast   (cl_axi_mstr_bus_4_q.wlast),
    .m_axi_wready  (cl_axi_mstr_bus_4_q.wready),
    .m_axi_bresp   (cl_axi_mstr_bus_4_q.bresp),
    .m_axi_bvalid  (cl_axi_mstr_bus_4_q.bvalid),
    .m_axi_bid     (cl_axi_mstr_bus_4_q.bid),
    .m_axi_bready  (cl_axi_mstr_bus_4_q.bready),
    .m_axi_arid    (cl_axi_mstr_bus_4_q.arid),
    .m_axi_araddr  (cl_axi_mstr_bus_4_q.araddr),
    .m_axi_arlen   (cl_axi_mstr_bus_4_q.arlen),
    .m_axi_arsize  (cl_axi_mstr_bus_4_q.arsize),
    .m_axi_arvalid (cl_axi_mstr_bus_4_q.arvalid),
    .m_axi_arready (cl_axi_mstr_bus_4_q.arready),
    .m_axi_rid     (cl_axi_mstr_bus_4_q.rid),
    .m_axi_rdata   (cl_axi_mstr_bus_4_q.rdata),
    .m_axi_rresp   (cl_axi_mstr_bus_4_q.rresp),
    .m_axi_rlast   (cl_axi_mstr_bus_4_q.rlast),
    .m_axi_rvalid  (cl_axi_mstr_bus_4_q.rvalid),
    .m_axi_rready  (cl_axi_mstr_bus_4_q.rready)
);
axi_register_slice MSTR_4_AXL_REG_SLC_2 (
    .aclk          (aclk),
    .aresetn       (aresetn),
    .s_axi_awid    (cl_axi_mstr_bus_4_q.awid),
    .s_axi_awaddr  (cl_axi_mstr_bus_4_q.awaddr),
    .s_axi_awlen   (cl_axi_mstr_bus_4_q.awlen),
    .s_axi_awvalid (cl_axi_mstr_bus_4_q.awvalid),
    .s_axi_awsize  (cl_axi_mstr_bus_4_q.awsize),
    .s_axi_awready (cl_axi_mstr_bus_4_q.awready),
    .s_axi_wdata   (cl_axi_mstr_bus_4_q.wdata),
    .s_axi_wstrb   (cl_axi_mstr_bus_4_q.wstrb),
    .s_axi_wlast   (cl_axi_mstr_bus_4_q.wlast),
    .s_axi_wvalid  (cl_axi_mstr_bus_4_q.wvalid),
    .s_axi_wready  (cl_axi_mstr_bus_4_q.wready),
    .s_axi_bid     (cl_axi_mstr_bus_4_q.bid),
    .s_axi_bresp   (cl_axi_mstr_bus_4_q.bresp),
    .s_axi_bvalid  (cl_axi_mstr_bus_4_q.bvalid),
    .s_axi_bready  (cl_axi_mstr_bus_4_q.bready),
    .s_axi_arid    (cl_axi_mstr_bus_4_q.arid),
    .s_axi_araddr  (cl_axi_mstr_bus_4_q.araddr),
    .s_axi_arlen   (cl_axi_mstr_bus_4_q.arlen),
    .s_axi_arvalid (cl_axi_mstr_bus_4_q.arvalid),
    .s_axi_arsize  (cl_axi_mstr_bus_4_q.arsize),
    .s_axi_arready (cl_axi_mstr_bus_4_q.arready),
    .s_axi_rid     (cl_axi_mstr_bus_4_q.rid),
    .s_axi_rdata   (cl_axi_mstr_bus_4_q.rdata),
    .s_axi_rresp   (cl_axi_mstr_bus_4_q.rresp),
    .s_axi_rlast   (cl_axi_mstr_bus_4_q.rlast),
    .s_axi_rvalid  (cl_axi_mstr_bus_4_q.rvalid),
    .s_axi_rready  (cl_axi_mstr_bus_4_q.rready),
    
    .m_axi_awid    (cl_axi_mstr_bus_4_q2.awid),
    .m_axi_awaddr  (cl_axi_mstr_bus_4_q2.awaddr),
    .m_axi_awlen   (cl_axi_mstr_bus_4_q2.awlen),
    .m_axi_awvalid (cl_axi_mstr_bus_4_q2.awvalid),
    .m_axi_awsize  (cl_axi_mstr_bus_4_q2.awsize),
    .m_axi_awready (cl_axi_mstr_bus_4_q2.awready),
    .m_axi_wdata   (cl_axi_mstr_bus_4_q2.wdata),
    .m_axi_wstrb   (cl_axi_mstr_bus_4_q2.wstrb),
    .m_axi_wvalid  (cl_axi_mstr_bus_4_q2.wvalid),
    .m_axi_wlast   (cl_axi_mstr_bus_4_q2.wlast),
    .m_axi_wready  (cl_axi_mstr_bus_4_q2.wready),
    .m_axi_bresp   (cl_axi_mstr_bus_4_q2.bresp),
    .m_axi_bvalid  (cl_axi_mstr_bus_4_q2.bvalid),
    .m_axi_bid     (cl_axi_mstr_bus_4_q2.bid),
    .m_axi_bready  (cl_axi_mstr_bus_4_q2.bready),
    .m_axi_arid    (cl_axi_mstr_bus_4_q2.arid),
    .m_axi_araddr  (cl_axi_mstr_bus_4_q2.araddr),
    .m_axi_arlen   (cl_axi_mstr_bus_4_q2.arlen),
    .m_axi_arsize  (cl_axi_mstr_bus_4_q2.arsize),
    .m_axi_arvalid (cl_axi_mstr_bus_4_q2.arvalid),
    .m_axi_arready (cl_axi_mstr_bus_4_q2.arready),
    .m_axi_rid     (cl_axi_mstr_bus_4_q2.rid),
    .m_axi_rdata   (cl_axi_mstr_bus_4_q2.rdata),
    .m_axi_rresp   (cl_axi_mstr_bus_4_q2.rresp),
    .m_axi_rlast   (cl_axi_mstr_bus_4_q2.rlast),
    .m_axi_rvalid  (cl_axi_mstr_bus_4_q2.rvalid),
    .m_axi_rready  (cl_axi_mstr_bus_4_q2.rready)
);


//----------------------------
// axi address translation modules
//----------------------------
axi_tlb #(
    .SR_ID(0)
) tlb1 (
    .clk(aclk),
    .rst(~aresetn),

    .virt_m(cl_axi_mstr_bus_1_q2),
    .phys_s(cl_axi_mstr_bus_1_t)
);
axi_tlb #(
    .SR_ID(1)
) tlb2 (
    .clk(aclk),
    .rst(~aresetn),

    .virt_m(cl_axi_mstr_bus_2_q2),
    .phys_s(cl_axi_mstr_bus_2_t)
);
axi_tlb #(
    .SR_ID(2)
) tlb3 (
    .clk(aclk),
    .rst(~aresetn),

    .virt_m(cl_axi_mstr_bus_3_q2),
    .phys_s(cl_axi_mstr_bus_3_t)
);
axi_tlb #(
    .SR_ID(3)
)  tlb4 (
    .clk(aclk),
    .rst(~aresetn),

    .virt_m(cl_axi_mstr_bus_4_q2),
    .phys_s(cl_axi_mstr_bus_4_t)
);


//----------------------------
// axi interconnect for DDR address decodes
//----------------------------
(* dont_touch = "true" *) cl_axi_interconnect AXI_CROSSBAR (
    .ACLK(aclk),
    .ARESETN(aresetn),

    .M00_AXI_araddr(lcl_cl_sh_ddra_q.araddr),
    .M00_AXI_arburst(),
    .M00_AXI_arcache(),
    .M00_AXI_arid(lcl_cl_sh_ddra_q.arid[8:0]),
    .M00_AXI_arlen(lcl_cl_sh_ddra_q.arlen),
    .M00_AXI_arlock(),
    .M00_AXI_arprot(),
    .M00_AXI_arqos(),
    .M00_AXI_arready(lcl_cl_sh_ddra_q.arready),
    .M00_AXI_arregion(),
    .M00_AXI_arsize(lcl_cl_sh_ddra_q.arsize),
    .M00_AXI_arvalid(lcl_cl_sh_ddra_q.arvalid),
    .M00_AXI_awaddr(lcl_cl_sh_ddra_q.awaddr),
    .M00_AXI_awburst(),
    .M00_AXI_awcache(),
    .M00_AXI_awid(lcl_cl_sh_ddra_q.awid[8:0]),
    .M00_AXI_awlen(lcl_cl_sh_ddra_q.awlen),
    .M00_AXI_awlock(),
    .M00_AXI_awprot(),
    .M00_AXI_awqos(),
    .M00_AXI_awready(lcl_cl_sh_ddra_q.awready),
    .M00_AXI_awregion(),
    .M00_AXI_awsize(lcl_cl_sh_ddra_q.awsize),
    .M00_AXI_awvalid(lcl_cl_sh_ddra_q.awvalid),
    .M00_AXI_bid(lcl_cl_sh_ddra_q.bid[8:0]),
    .M00_AXI_bready(lcl_cl_sh_ddra_q.bready),
    .M00_AXI_bresp(lcl_cl_sh_ddra_q.bresp),
    .M00_AXI_bvalid(lcl_cl_sh_ddra_q.bvalid),
    .M00_AXI_rdata(lcl_cl_sh_ddra_q.rdata),
    .M00_AXI_rid(lcl_cl_sh_ddra_q.rid[8:0]),
    .M00_AXI_rlast(lcl_cl_sh_ddra_q.rlast),
    .M00_AXI_rready(lcl_cl_sh_ddra_q.rready),
    .M00_AXI_rresp(lcl_cl_sh_ddra_q.rresp),
    .M00_AXI_rvalid(lcl_cl_sh_ddra_q.rvalid),
    .M00_AXI_wdata(lcl_cl_sh_ddra_q.wdata),
    .M00_AXI_wlast(lcl_cl_sh_ddra_q.wlast),
    .M00_AXI_wready(lcl_cl_sh_ddra_q.wready),
    .M00_AXI_wstrb(lcl_cl_sh_ddra_q.wstrb),
    .M00_AXI_wvalid(lcl_cl_sh_ddra_q.wvalid),

    .M01_AXI_araddr(lcl_cl_sh_ddrb_q.araddr),
    .M01_AXI_arburst(),
    .M01_AXI_arcache(),
    .M01_AXI_arid(lcl_cl_sh_ddrb_q.arid[8:0]),
    .M01_AXI_arlen(lcl_cl_sh_ddrb_q.arlen),
    .M01_AXI_arlock(),
    .M01_AXI_arprot(),
    .M01_AXI_arqos(),
    .M01_AXI_arready(lcl_cl_sh_ddrb_q.arready),
    .M01_AXI_arregion(),
    .M01_AXI_arsize(lcl_cl_sh_ddrb_q.arsize),
    .M01_AXI_arvalid(lcl_cl_sh_ddrb_q.arvalid),
    .M01_AXI_awaddr(lcl_cl_sh_ddrb_q.awaddr),
    .M01_AXI_awburst(),
    .M01_AXI_awcache(),
    .M01_AXI_awid(lcl_cl_sh_ddrb_q.awid[8:0]),
    .M01_AXI_awlen(lcl_cl_sh_ddrb_q.awlen),
    .M01_AXI_awlock(),
    .M01_AXI_awprot(),
    .M01_AXI_awqos(),
    .M01_AXI_awready(lcl_cl_sh_ddrb_q.awready),
    .M01_AXI_awregion(),
    .M01_AXI_awsize(lcl_cl_sh_ddrb_q.awsize),
    .M01_AXI_awvalid(lcl_cl_sh_ddrb_q.awvalid),
    .M01_AXI_bid(lcl_cl_sh_ddrb_q.bid[8:0]),
    .M01_AXI_bready(lcl_cl_sh_ddrb_q.bready),
    .M01_AXI_bresp(lcl_cl_sh_ddrb_q.bresp),
    .M01_AXI_bvalid(lcl_cl_sh_ddrb_q.bvalid),
    .M01_AXI_rdata(lcl_cl_sh_ddrb_q.rdata),
    .M01_AXI_rid(lcl_cl_sh_ddrb_q.rid[8:0]),
    .M01_AXI_rlast(lcl_cl_sh_ddrb_q.rlast),
    .M01_AXI_rready(lcl_cl_sh_ddrb_q.rready),
    .M01_AXI_rresp(lcl_cl_sh_ddrb_q.rresp),
    .M01_AXI_rvalid(lcl_cl_sh_ddrb_q.rvalid),
    .M01_AXI_wdata(lcl_cl_sh_ddrb_q.wdata),
    .M01_AXI_wlast(lcl_cl_sh_ddrb_q.wlast),
    .M01_AXI_wready(lcl_cl_sh_ddrb_q.wready),
    .M01_AXI_wstrb(lcl_cl_sh_ddrb_q.wstrb),
    .M01_AXI_wvalid(lcl_cl_sh_ddrb_q.wvalid),

    .M02_AXI_araddr(cl_sh_ddr_q.araddr),
    .M02_AXI_arburst(),
    .M02_AXI_arcache(),
    .M02_AXI_arid(cl_sh_ddr_q.arid[8:0]),
    .M02_AXI_arlen(cl_sh_ddr_q.arlen),
    .M02_AXI_arlock(),
    .M02_AXI_arprot(),
    .M02_AXI_arqos(),
    .M02_AXI_arready(cl_sh_ddr_q.arready),
    .M02_AXI_arregion(),
    .M02_AXI_arsize(cl_sh_ddr_q.arsize),
    .M02_AXI_arvalid(cl_sh_ddr_q.arvalid),
    .M02_AXI_awaddr(cl_sh_ddr_q.awaddr),
    .M02_AXI_awburst(),
    .M02_AXI_awcache(),
    .M02_AXI_awid(cl_sh_ddr_q.awid[8:0]),
    .M02_AXI_awlen(cl_sh_ddr_q.awlen),
    .M02_AXI_awlock(),
    .M02_AXI_awprot(),
    .M02_AXI_awqos(),
    .M02_AXI_awready(cl_sh_ddr_q.awready),
    .M02_AXI_awregion(),
    .M02_AXI_awsize(cl_sh_ddr_q.awsize),
    .M02_AXI_awvalid(cl_sh_ddr_q.awvalid),
    .M02_AXI_bid(cl_sh_ddr_q.bid[8:0]),
    .M02_AXI_bready(cl_sh_ddr_q.bready),
    .M02_AXI_bresp(cl_sh_ddr_q.bresp),
    .M02_AXI_bvalid(cl_sh_ddr_q.bvalid),
    .M02_AXI_rdata(cl_sh_ddr_q.rdata),
    .M02_AXI_rid(cl_sh_ddr_q.rid[8:0]),
    .M02_AXI_rlast(cl_sh_ddr_q.rlast),
    .M02_AXI_rready(cl_sh_ddr_q.rready),
    .M02_AXI_rresp(cl_sh_ddr_q.rresp),
    .M02_AXI_rvalid(cl_sh_ddr_q.rvalid),
    .M02_AXI_wdata(cl_sh_ddr_q.wdata),
    .M02_AXI_wlast(cl_sh_ddr_q.wlast),
    .M02_AXI_wready(cl_sh_ddr_q.wready),
    .M02_AXI_wstrb(cl_sh_ddr_q.wstrb),
    .M02_AXI_wvalid(cl_sh_ddr_q.wvalid),

    .M03_AXI_araddr(lcl_cl_sh_ddrd_q.araddr),
    .M03_AXI_arburst(),
    .M03_AXI_arcache(),
    .M03_AXI_arid(lcl_cl_sh_ddrd_q.arid[8:0]),
    .M03_AXI_arlen(lcl_cl_sh_ddrd_q.arlen),
    .M03_AXI_arlock(),
    .M03_AXI_arprot(),
    .M03_AXI_arqos(),
    .M03_AXI_arready(lcl_cl_sh_ddrd_q.arready),
    .M03_AXI_arregion(),
    .M03_AXI_arsize(lcl_cl_sh_ddrd_q.arsize),
    .M03_AXI_arvalid(lcl_cl_sh_ddrd_q.arvalid),
    .M03_AXI_awaddr(lcl_cl_sh_ddrd_q.awaddr),
    .M03_AXI_awburst(),
    .M03_AXI_awcache(),
    .M03_AXI_awid(lcl_cl_sh_ddrd_q.awid[8:0]),
    .M03_AXI_awlen(lcl_cl_sh_ddrd_q.awlen),
    .M03_AXI_awlock(),
    .M03_AXI_awprot(),
    .M03_AXI_awqos(),
    .M03_AXI_awready(lcl_cl_sh_ddrd_q.awready),
    .M03_AXI_awregion(),
    .M03_AXI_awsize(lcl_cl_sh_ddrd_q.awsize),
    .M03_AXI_awvalid(lcl_cl_sh_ddrd_q.awvalid),
    .M03_AXI_bid(lcl_cl_sh_ddrd_q.bid[8:0]),
    .M03_AXI_bready(lcl_cl_sh_ddrd_q.bready),
    .M03_AXI_bresp(lcl_cl_sh_ddrd_q.bresp),
    .M03_AXI_bvalid(lcl_cl_sh_ddrd_q.bvalid),
    .M03_AXI_rdata(lcl_cl_sh_ddrd_q.rdata),
    .M03_AXI_rid(lcl_cl_sh_ddrd_q.rid[8:0]),
    .M03_AXI_rlast(lcl_cl_sh_ddrd_q.rlast),
    .M03_AXI_rready(lcl_cl_sh_ddrd_q.rready),
    .M03_AXI_rresp(lcl_cl_sh_ddrd_q.rresp),
    .M03_AXI_rvalid(lcl_cl_sh_ddrd_q.rvalid),
    .M03_AXI_wdata(lcl_cl_sh_ddrd_q.wdata),
    .M03_AXI_wlast(lcl_cl_sh_ddrd_q.wlast),
    .M03_AXI_wready(lcl_cl_sh_ddrd_q.wready),
    .M03_AXI_wstrb(lcl_cl_sh_ddrd_q.wstrb),
    .M03_AXI_wvalid(lcl_cl_sh_ddrd_q.wvalid),

    .S00_AXI_araddr({sh_cl_dma_pcis_q.araddr[63:37], 1'b0, sh_cl_dma_pcis_q.araddr[35:0]}),
    .S00_AXI_arburst(2'b1),
    .S00_AXI_arcache(4'b11),
    .S00_AXI_arid(sh_cl_dma_pcis_q.arid[5:0]),
    .S00_AXI_arlen(sh_cl_dma_pcis_q.arlen),
    .S00_AXI_arlock(1'b0),
    .S00_AXI_arprot(3'b10),
    .S00_AXI_arqos(4'b0),
    .S00_AXI_arready(sh_cl_dma_pcis_q.arready),
    .S00_AXI_arregion(4'b0),
    .S00_AXI_arsize(sh_cl_dma_pcis_q.arsize),
    .S00_AXI_arvalid(sh_cl_dma_pcis_q.arvalid),
    .S00_AXI_awaddr({sh_cl_dma_pcis_q.awaddr[63:37], 1'b0, sh_cl_dma_pcis_q.awaddr[35:0]}),
    .S00_AXI_awburst(2'b1),
    .S00_AXI_awcache(4'b11),
    .S00_AXI_awid(sh_cl_dma_pcis_q.awid[5:0]),
    .S00_AXI_awlen(sh_cl_dma_pcis_q.awlen),
    .S00_AXI_awlock(1'b0),
    .S00_AXI_awprot(3'b10),
    .S00_AXI_awqos(4'b0),
    .S00_AXI_awready(sh_cl_dma_pcis_q.awready),
    .S00_AXI_awregion(4'b0),
    .S00_AXI_awsize(sh_cl_dma_pcis_q.awsize),
    .S00_AXI_awvalid(sh_cl_dma_pcis_q.awvalid),
    .S00_AXI_bid(sh_cl_dma_pcis_q.bid[5:0]),
    .S00_AXI_bready(sh_cl_dma_pcis_q.bready),
    .S00_AXI_bresp(sh_cl_dma_pcis_q.bresp),
    .S00_AXI_bvalid(sh_cl_dma_pcis_q.bvalid),
    .S00_AXI_rdata(sh_cl_dma_pcis_q.rdata),
    .S00_AXI_rid(sh_cl_dma_pcis_q.rid[5:0]),
    .S00_AXI_rlast(sh_cl_dma_pcis_q.rlast),
    .S00_AXI_rready(sh_cl_dma_pcis_q.rready),
    .S00_AXI_rresp(sh_cl_dma_pcis_q.rresp),
    .S00_AXI_rvalid(sh_cl_dma_pcis_q.rvalid),
    .S00_AXI_wdata(sh_cl_dma_pcis_q.wdata),
    .S00_AXI_wlast(sh_cl_dma_pcis_q.wlast),
    .S00_AXI_wready(sh_cl_dma_pcis_q.wready),
    .S00_AXI_wstrb(sh_cl_dma_pcis_q.wstrb),
    .S00_AXI_wvalid(sh_cl_dma_pcis_q.wvalid),

    .S01_AXI_araddr({cl_axi_mstr_bus_1_t.araddr}),
    .S01_AXI_arburst(2'b1),
    .S01_AXI_arcache(4'b11),
    .S01_AXI_arid(cl_axi_mstr_bus_1_t.arid[6:0]),
    .S01_AXI_arlen(cl_axi_mstr_bus_1_t.arlen),
    .S01_AXI_arlock(1'b0),
    .S01_AXI_arprot(3'b10),
    .S01_AXI_arqos(4'b0),
    .S01_AXI_arready(cl_axi_mstr_bus_1_t.arready),
    .S01_AXI_arregion(4'b0),
    .S01_AXI_arsize(cl_axi_mstr_bus_1_t.arsize),
    .S01_AXI_arvalid(cl_axi_mstr_bus_1_t.arvalid),
    .S01_AXI_awaddr({cl_axi_mstr_bus_1_t.awaddr}),
    .S01_AXI_awburst(2'b1),
    .S01_AXI_awcache(4'b11),
    .S01_AXI_awid(cl_axi_mstr_bus_1_t.awid[6:0]),
    .S01_AXI_awlen(cl_axi_mstr_bus_1_t.awlen),
    .S01_AXI_awlock(1'b0),
    .S01_AXI_awprot(3'b10),
    .S01_AXI_awqos(4'b0),
    .S01_AXI_awready(cl_axi_mstr_bus_1_t.awready),
    .S01_AXI_awregion(4'b0),
    .S01_AXI_awsize(cl_axi_mstr_bus_1_t.awsize),
    .S01_AXI_awvalid(cl_axi_mstr_bus_1_t.awvalid),
    .S01_AXI_bid(cl_axi_mstr_bus_1_t.bid[6:0]),
    .S01_AXI_bready(cl_axi_mstr_bus_1_t.bready),
    .S01_AXI_bresp(cl_axi_mstr_bus_1_t.bresp),
    .S01_AXI_bvalid(cl_axi_mstr_bus_1_t.bvalid),
    .S01_AXI_rdata(cl_axi_mstr_bus_1_t.rdata),
    .S01_AXI_rid(cl_axi_mstr_bus_1_t.rid[6:0]),
    .S01_AXI_rlast(cl_axi_mstr_bus_1_t.rlast),
    .S01_AXI_rready(cl_axi_mstr_bus_1_t.rready),
    .S01_AXI_rresp(cl_axi_mstr_bus_1_t.rresp),
    .S01_AXI_rvalid(cl_axi_mstr_bus_1_t.rvalid),
    .S01_AXI_wdata(cl_axi_mstr_bus_1_t.wdata),
    .S01_AXI_wlast(cl_axi_mstr_bus_1_t.wlast),
    .S01_AXI_wready(cl_axi_mstr_bus_1_t.wready),
    .S01_AXI_wstrb(cl_axi_mstr_bus_1_t.wstrb),
    .S01_AXI_wvalid(cl_axi_mstr_bus_1_t.wvalid),

    .S02_AXI_araddr({cl_axi_mstr_bus_2_t.araddr}),
    .S02_AXI_arburst(2'b1),
    .S02_AXI_arcache(4'b11),
    .S02_AXI_arid(cl_axi_mstr_bus_2_t.arid[6:0]),
    .S02_AXI_arlen(cl_axi_mstr_bus_2_t.arlen),
    .S02_AXI_arlock(1'b0),
    .S02_AXI_arprot(3'b10),
    .S02_AXI_arqos(4'b0),
    .S02_AXI_arready(cl_axi_mstr_bus_2_t.arready),
    .S02_AXI_arregion(4'b0),
    .S02_AXI_arsize(cl_axi_mstr_bus_2_t.arsize),
    .S02_AXI_arvalid(cl_axi_mstr_bus_2_t.arvalid),
    .S02_AXI_awaddr({cl_axi_mstr_bus_2_t.awaddr}),
    .S02_AXI_awburst(2'b1),
    .S02_AXI_awcache(4'b11),
    .S02_AXI_awid(cl_axi_mstr_bus_2_t.awid[6:0]),
    .S02_AXI_awlen(cl_axi_mstr_bus_2_t.awlen),
    .S02_AXI_awlock(1'b0),
    .S02_AXI_awprot(3'b10),
    .S02_AXI_awqos(4'b0),
    .S02_AXI_awready(cl_axi_mstr_bus_2_t.awready),
    .S02_AXI_awregion(4'b0),
    .S02_AXI_awsize(cl_axi_mstr_bus_2_t.awsize),
    .S02_AXI_awvalid(cl_axi_mstr_bus_2_t.awvalid),
    .S02_AXI_bid(cl_axi_mstr_bus_2_t.bid[6:0]),
    .S02_AXI_bready(cl_axi_mstr_bus_2_t.bready),
    .S02_AXI_bresp(cl_axi_mstr_bus_2_t.bresp),
    .S02_AXI_bvalid(cl_axi_mstr_bus_2_t.bvalid),
    .S02_AXI_rdata(cl_axi_mstr_bus_2_t.rdata),
    .S02_AXI_rid(cl_axi_mstr_bus_2_t.rid[6:0]),
    .S02_AXI_rlast(cl_axi_mstr_bus_2_t.rlast),
    .S02_AXI_rready(cl_axi_mstr_bus_2_t.rready),
    .S02_AXI_rresp(cl_axi_mstr_bus_2_t.rresp),
    .S02_AXI_rvalid(cl_axi_mstr_bus_2_t.rvalid),
    .S02_AXI_wdata(cl_axi_mstr_bus_2_t.wdata),
    .S02_AXI_wlast(cl_axi_mstr_bus_2_t.wlast),
    .S02_AXI_wready(cl_axi_mstr_bus_2_t.wready),
    .S02_AXI_wstrb(cl_axi_mstr_bus_2_t.wstrb),
    .S02_AXI_wvalid(cl_axi_mstr_bus_2_t.wvalid),

    .S03_AXI_araddr({cl_axi_mstr_bus_3_t.araddr}),
    .S03_AXI_arburst(2'b1),
    .S03_AXI_arcache(4'b11),
    .S03_AXI_arid(cl_axi_mstr_bus_3_t.arid[6:0]),
    .S03_AXI_arlen(cl_axi_mstr_bus_3_t.arlen),
    .S03_AXI_arlock(1'b0),
    .S03_AXI_arprot(3'b10),
    .S03_AXI_arqos(4'b0),
    .S03_AXI_arready(cl_axi_mstr_bus_3_t.arready),
    .S03_AXI_arregion(4'b0),
    .S03_AXI_arsize(cl_axi_mstr_bus_3_t.arsize),
    .S03_AXI_arvalid(cl_axi_mstr_bus_3_t.arvalid),
    .S03_AXI_awaddr({cl_axi_mstr_bus_3_t.awaddr}),
    .S03_AXI_awburst(2'b1),
    .S03_AXI_awcache(4'b11),
    .S03_AXI_awid(cl_axi_mstr_bus_3_t.awid[6:0]),
    .S03_AXI_awlen(cl_axi_mstr_bus_3_t.awlen),
    .S03_AXI_awlock(1'b0),
    .S03_AXI_awprot(3'b10),
    .S03_AXI_awqos(4'b0),
    .S03_AXI_awready(cl_axi_mstr_bus_3_t.awready),
    .S03_AXI_awregion(4'b0),
    .S03_AXI_awsize(cl_axi_mstr_bus_3_t.awsize),
    .S03_AXI_awvalid(cl_axi_mstr_bus_3_t.awvalid),
    .S03_AXI_bid(cl_axi_mstr_bus_3_t.bid[6:0]),
    .S03_AXI_bready(cl_axi_mstr_bus_3_t.bready),
    .S03_AXI_bresp(cl_axi_mstr_bus_3_t.bresp),
    .S03_AXI_bvalid(cl_axi_mstr_bus_3_t.bvalid),
    .S03_AXI_rdata(cl_axi_mstr_bus_3_t.rdata),
    .S03_AXI_rid(cl_axi_mstr_bus_3_t.rid[6:0]),
    .S03_AXI_rlast(cl_axi_mstr_bus_3_t.rlast),
    .S03_AXI_rready(cl_axi_mstr_bus_3_t.rready),
    .S03_AXI_rresp(cl_axi_mstr_bus_3_t.rresp),
    .S03_AXI_rvalid(cl_axi_mstr_bus_3_t.rvalid),
    .S03_AXI_wdata(cl_axi_mstr_bus_3_t.wdata),
    .S03_AXI_wlast(cl_axi_mstr_bus_3_t.wlast),
    .S03_AXI_wready(cl_axi_mstr_bus_3_t.wready),
    .S03_AXI_wstrb(cl_axi_mstr_bus_3_t.wstrb),
    .S03_AXI_wvalid(cl_axi_mstr_bus_3_t.wvalid),

    .S04_AXI_araddr({cl_axi_mstr_bus_4_t.araddr}),
    .S04_AXI_arburst(2'b1),
    .S04_AXI_arcache(4'b11),
    .S04_AXI_arid(cl_axi_mstr_bus_4_t.arid[6:0]),
    .S04_AXI_arlen(cl_axi_mstr_bus_4_t.arlen),
    .S04_AXI_arlock(1'b0),
    .S04_AXI_arprot(3'b10),
    .S04_AXI_arqos(4'b0),
    .S04_AXI_arready(cl_axi_mstr_bus_4_t.arready),
    .S04_AXI_arregion(4'b0),
    .S04_AXI_arsize(cl_axi_mstr_bus_4_t.arsize),
    .S04_AXI_arvalid(cl_axi_mstr_bus_4_t.arvalid),
    .S04_AXI_awaddr({cl_axi_mstr_bus_4_t.awaddr}),
    .S04_AXI_awburst(2'b1),
    .S04_AXI_awcache(4'b11),
    .S04_AXI_awid(cl_axi_mstr_bus_4_t.awid[6:0]),
    .S04_AXI_awlen(cl_axi_mstr_bus_4_t.awlen),
    .S04_AXI_awlock(1'b0),
    .S04_AXI_awprot(3'b10),
    .S04_AXI_awqos(4'b0),
    .S04_AXI_awready(cl_axi_mstr_bus_4_t.awready),
    .S04_AXI_awregion(4'b0),
    .S04_AXI_awsize(cl_axi_mstr_bus_4_t.awsize),
    .S04_AXI_awvalid(cl_axi_mstr_bus_4_t.awvalid),
    .S04_AXI_bid(cl_axi_mstr_bus_4_t.bid[6:0]),
    .S04_AXI_bready(cl_axi_mstr_bus_4_t.bready),
    .S04_AXI_bresp(cl_axi_mstr_bus_4_t.bresp),
    .S04_AXI_bvalid(cl_axi_mstr_bus_4_t.bvalid),
    .S04_AXI_rdata(cl_axi_mstr_bus_4_t.rdata),
    .S04_AXI_rid(cl_axi_mstr_bus_4_t.rid[6:0]),
    .S04_AXI_rlast(cl_axi_mstr_bus_4_t.rlast),
    .S04_AXI_rready(cl_axi_mstr_bus_4_t.rready),
    .S04_AXI_rresp(cl_axi_mstr_bus_4_t.rresp),
    .S04_AXI_rvalid(cl_axi_mstr_bus_4_t.rvalid),
    .S04_AXI_wdata(cl_axi_mstr_bus_4_t.wdata),
    .S04_AXI_wlast(cl_axi_mstr_bus_4_t.wlast),
    .S04_AXI_wready(cl_axi_mstr_bus_4_t.wready),
    .S04_AXI_wstrb(cl_axi_mstr_bus_4_t.wstrb),
    .S04_AXI_wvalid(cl_axi_mstr_bus_4_t.wvalid)
);

//----------------------------
// flop the output of interconnect for DDRC
//----------------------------
src_register_slice DDR_C_TST_AXI4_REG_SLC (
    .aclk           (aclk),
    .aresetn        (aresetn),

    .s_axi_awid     (cl_sh_ddr_q.awid),
    .s_axi_awaddr   ({cl_sh_ddr_q.awaddr[63:36], 2'b0, cl_sh_ddr_q.awaddr[33:0]}),
    .s_axi_awlen    (cl_sh_ddr_q.awlen),
    .s_axi_awsize   (cl_sh_ddr_q.awsize),
    .s_axi_awvalid  (cl_sh_ddr_q.awvalid),
    .s_axi_awready  (cl_sh_ddr_q.awready),
    .s_axi_wdata    (cl_sh_ddr_q.wdata),
    .s_axi_wstrb    (cl_sh_ddr_q.wstrb),
    .s_axi_wlast    (cl_sh_ddr_q.wlast),
    .s_axi_wvalid   (cl_sh_ddr_q.wvalid),
    .s_axi_wready   (cl_sh_ddr_q.wready),
    .s_axi_bid      (cl_sh_ddr_q.bid),
    .s_axi_bresp    (cl_sh_ddr_q.bresp),
    .s_axi_bvalid   (cl_sh_ddr_q.bvalid),
    .s_axi_bready   (cl_sh_ddr_q.bready),
    .s_axi_arid     (cl_sh_ddr_q.arid),
    .s_axi_araddr   ({cl_sh_ddr_q.araddr[63:36], 2'b0, cl_sh_ddr_q.araddr[33:0]}),
    .s_axi_arlen    (cl_sh_ddr_q.arlen),
    .s_axi_arsize   (cl_sh_ddr_q.arsize),
    .s_axi_arvalid  (cl_sh_ddr_q.arvalid),
    .s_axi_arready  (cl_sh_ddr_q.arready),
    .s_axi_rid      (cl_sh_ddr_q.rid),
    .s_axi_rdata    (cl_sh_ddr_q.rdata),
    .s_axi_rresp    (cl_sh_ddr_q.rresp),
    .s_axi_rlast    (cl_sh_ddr_q.rlast),
    .s_axi_rvalid   (cl_sh_ddr_q.rvalid),
    .s_axi_rready   (cl_sh_ddr_q.rready),
    
    .m_axi_awid     (cl_sh_ddr_q2.awid),
    .m_axi_awaddr   (cl_sh_ddr_q2.awaddr),
    .m_axi_awlen    (cl_sh_ddr_q2.awlen),
    .m_axi_awsize   (cl_sh_ddr_q2.awsize),
    .m_axi_awvalid  (cl_sh_ddr_q2.awvalid),
    .m_axi_awready  (cl_sh_ddr_q2.awready),
    .m_axi_wdata    (cl_sh_ddr_q2.wdata),
    .m_axi_wstrb    (cl_sh_ddr_q2.wstrb),
    .m_axi_wlast    (cl_sh_ddr_q2.wlast),
    .m_axi_wvalid   (cl_sh_ddr_q2.wvalid),
    .m_axi_wready   (cl_sh_ddr_q2.wready),
    .m_axi_bid      (cl_sh_ddr_q2.bid),
    .m_axi_bresp    (cl_sh_ddr_q2.bresp),
    .m_axi_bvalid   (cl_sh_ddr_q2.bvalid),
    .m_axi_bready   (cl_sh_ddr_q2.bready),
    .m_axi_arid     (cl_sh_ddr_q2.arid),
    .m_axi_araddr   (cl_sh_ddr_q2.araddr),
    .m_axi_arlen    (cl_sh_ddr_q2.arlen),
    .m_axi_arsize   (cl_sh_ddr_q2.arsize),
    .m_axi_arvalid  (cl_sh_ddr_q2.arvalid),
    .m_axi_arready  (cl_sh_ddr_q2.arready),
    .m_axi_rid      (cl_sh_ddr_q2.rid),
    .m_axi_rdata    (cl_sh_ddr_q2.rdata),
    .m_axi_rresp    (cl_sh_ddr_q2.rresp),
    .m_axi_rlast    (cl_sh_ddr_q2.rlast),
    .m_axi_rvalid   (cl_sh_ddr_q2.rvalid),
    .m_axi_rready   (cl_sh_ddr_q2.rready)
);

dest_register_slice DDR_C_TST_AXI4_REG_SLC_1 (
    .aclk           (aclk),
    .aresetn        (aresetn),
  
    .s_axi_awid     (cl_sh_ddr_q2.awid),
    .s_axi_awaddr   (cl_sh_ddr_q2.awaddr),
    .s_axi_awlen    (cl_sh_ddr_q2.awlen),
    .s_axi_awsize   (cl_sh_ddr_q2.awsize),
    .s_axi_awvalid  (cl_sh_ddr_q2.awvalid),
    .s_axi_awready  (cl_sh_ddr_q2.awready),
    .s_axi_wdata    (cl_sh_ddr_q2.wdata),
    .s_axi_wstrb    (cl_sh_ddr_q2.wstrb),
    .s_axi_wlast    (cl_sh_ddr_q2.wlast),
    .s_axi_wvalid   (cl_sh_ddr_q2.wvalid),
    .s_axi_wready   (cl_sh_ddr_q2.wready),
    .s_axi_bid      (cl_sh_ddr_q2.bid),
    .s_axi_bresp    (cl_sh_ddr_q2.bresp),
    .s_axi_bvalid   (cl_sh_ddr_q2.bvalid),
    .s_axi_bready   (cl_sh_ddr_q2.bready),
    .s_axi_arid     (cl_sh_ddr_q2.arid),
    .s_axi_araddr   (cl_sh_ddr_q2.araddr),
    .s_axi_arlen    (cl_sh_ddr_q2.arlen),
    .s_axi_arsize   (cl_sh_ddr_q2.arsize),
    .s_axi_arvalid  (cl_sh_ddr_q2.arvalid),
    .s_axi_arready  (cl_sh_ddr_q2.arready),
    .s_axi_rid      (cl_sh_ddr_q2.rid),
    .s_axi_rdata    (cl_sh_ddr_q2.rdata),
    .s_axi_rresp    (cl_sh_ddr_q2.rresp),
    .s_axi_rlast    (cl_sh_ddr_q2.rlast),
    .s_axi_rvalid   (cl_sh_ddr_q2.rvalid),
    .s_axi_rready   (cl_sh_ddr_q2.rready),
  
    .m_axi_awid     (cl_sh_ddr_bus.awid),
    .m_axi_awaddr   (cl_sh_ddr_bus.awaddr),
    .m_axi_awlen    (cl_sh_ddr_bus.awlen),
    .m_axi_awsize   (cl_sh_ddr_bus.awsize),
    .m_axi_awvalid  (cl_sh_ddr_bus.awvalid),
    .m_axi_awready  (cl_sh_ddr_bus.awready),
    .m_axi_wdata    (cl_sh_ddr_bus.wdata),
    .m_axi_wstrb    (cl_sh_ddr_bus.wstrb),
    .m_axi_wlast    (cl_sh_ddr_bus.wlast),
    .m_axi_wvalid   (cl_sh_ddr_bus.wvalid),
    .m_axi_wready   (cl_sh_ddr_bus.wready),
    .m_axi_bid      (cl_sh_ddr_bus.bid),
    .m_axi_bresp    (cl_sh_ddr_bus.bresp),
    .m_axi_bvalid   (cl_sh_ddr_bus.bvalid),
    .m_axi_bready   (cl_sh_ddr_bus.bready),
    .m_axi_arid     (cl_sh_ddr_bus.arid),
    .m_axi_araddr   (cl_sh_ddr_bus.araddr),
    .m_axi_arlen    (cl_sh_ddr_bus.arlen),
    .m_axi_arsize   (cl_sh_ddr_bus.arsize),
    .m_axi_arvalid  (cl_sh_ddr_bus.arvalid),
    .m_axi_arready  (cl_sh_ddr_bus.arready),
    .m_axi_rid      (cl_sh_ddr_bus.rid),
    .m_axi_rdata    (cl_sh_ddr_bus.rdata),
    .m_axi_rresp    (cl_sh_ddr_bus.rresp),
    .m_axi_rlast    (cl_sh_ddr_bus.rlast),
    .m_axi_rvalid   (cl_sh_ddr_bus.rvalid),
    .m_axi_rready   (cl_sh_ddr_bus.rready)
);


//----------------------------
// flop the output of interconnect for DDRA
// back to back for SLR crossing
//----------------------------
//back to back register slices for SLR crossing
src_register_slice DDR_A_TST_AXI4_REG_SLC_1 (
    .aclk           (aclk),
    .aresetn        (aresetn),
    .s_axi_awid     (lcl_cl_sh_ddra_q.awid),
    .s_axi_awaddr   ({lcl_cl_sh_ddra_q.awaddr[63:36], 2'b0, lcl_cl_sh_ddra_q.awaddr[33:0]}),
    .s_axi_awlen    (lcl_cl_sh_ddra_q.awlen),
    .s_axi_awsize   (lcl_cl_sh_ddra_q.awsize),
    .s_axi_awburst  (2'b1),
    .s_axi_awlock   (1'b0),
    .s_axi_awcache  (4'b11),
    .s_axi_awprot   (3'b10),
    .s_axi_awregion (4'b0),
    .s_axi_awqos    (4'b0),
    .s_axi_awvalid  (lcl_cl_sh_ddra_q.awvalid),
    .s_axi_awready  (lcl_cl_sh_ddra_q.awready),
    .s_axi_wdata    (lcl_cl_sh_ddra_q.wdata),
    .s_axi_wstrb    (lcl_cl_sh_ddra_q.wstrb),
    .s_axi_wlast    (lcl_cl_sh_ddra_q.wlast),
    .s_axi_wvalid   (lcl_cl_sh_ddra_q.wvalid),
    .s_axi_wready   (lcl_cl_sh_ddra_q.wready),
    .s_axi_bid      (lcl_cl_sh_ddra_q.bid),
    .s_axi_bresp    (lcl_cl_sh_ddra_q.bresp),
    .s_axi_bvalid   (lcl_cl_sh_ddra_q.bvalid),
    .s_axi_bready   (lcl_cl_sh_ddra_q.bready),
    .s_axi_arid     (lcl_cl_sh_ddra_q.arid),
    .s_axi_araddr   ({lcl_cl_sh_ddra_q.araddr[63:36], 2'b0, lcl_cl_sh_ddra_q.araddr[33:0]}),
    .s_axi_arlen    (lcl_cl_sh_ddra_q.arlen),
    .s_axi_arsize   (lcl_cl_sh_ddra_q.arsize),
    .s_axi_arburst  (2'b1),
    .s_axi_arlock   (1'b0),
    .s_axi_arcache  (4'b11),
    .s_axi_arprot   (3'b10),
    .s_axi_arregion (4'b0),
    .s_axi_arqos    (4'b0),
    .s_axi_arvalid  (lcl_cl_sh_ddra_q.arvalid),
    .s_axi_arready  (lcl_cl_sh_ddra_q.arready),
    .s_axi_rid      (lcl_cl_sh_ddra_q.rid),
    .s_axi_rdata    (lcl_cl_sh_ddra_q.rdata),
    .s_axi_rresp    (lcl_cl_sh_ddra_q.rresp),
    .s_axi_rlast    (lcl_cl_sh_ddra_q.rlast),
    .s_axi_rvalid   (lcl_cl_sh_ddra_q.rvalid),
    .s_axi_rready   (lcl_cl_sh_ddra_q.rready),
    
    .m_axi_awid     (lcl_cl_sh_ddra_q2.awid),
    .m_axi_awaddr   (lcl_cl_sh_ddra_q2.awaddr),
    .m_axi_awlen    (lcl_cl_sh_ddra_q2.awlen),
    .m_axi_awsize   (lcl_cl_sh_ddra_q2.awsize),
    .m_axi_awburst  (),
    .m_axi_awlock   (),
    .m_axi_awcache  (),
    .m_axi_awprot   (),
    .m_axi_awregion (),
    .m_axi_awqos    (),
    .m_axi_awvalid  (lcl_cl_sh_ddra_q2.awvalid),
    .m_axi_awready  (lcl_cl_sh_ddra_q2.awready),
    .m_axi_wdata    (lcl_cl_sh_ddra_q2.wdata),
    .m_axi_wstrb    (lcl_cl_sh_ddra_q2.wstrb),
    .m_axi_wlast    (lcl_cl_sh_ddra_q2.wlast),
    .m_axi_wvalid   (lcl_cl_sh_ddra_q2.wvalid),
    .m_axi_wready   (lcl_cl_sh_ddra_q2.wready),
    .m_axi_bid      (lcl_cl_sh_ddra_q2.bid),
    .m_axi_bresp    (lcl_cl_sh_ddra_q2.bresp),
    .m_axi_bvalid   (lcl_cl_sh_ddra_q2.bvalid),
    .m_axi_bready   (lcl_cl_sh_ddra_q2.bready),
    .m_axi_arid     (lcl_cl_sh_ddra_q2.arid),
    .m_axi_araddr   (lcl_cl_sh_ddra_q2.araddr),
    .m_axi_arlen    (lcl_cl_sh_ddra_q2.arlen),
    .m_axi_arsize   (lcl_cl_sh_ddra_q2.arsize),
    .m_axi_arburst  (),
    .m_axi_arlock   (),
    .m_axi_arcache  (),
    .m_axi_arprot   (),
    .m_axi_arregion (),
    .m_axi_arqos    (),
    .m_axi_arvalid  (lcl_cl_sh_ddra_q2.arvalid),
    .m_axi_arready  (lcl_cl_sh_ddra_q2.arready),
    .m_axi_rid      (lcl_cl_sh_ddra_q2.rid),
    .m_axi_rdata    (lcl_cl_sh_ddra_q2.rdata),
    .m_axi_rresp    (lcl_cl_sh_ddra_q2.rresp),
    .m_axi_rlast    (lcl_cl_sh_ddra_q2.rlast),
    .m_axi_rvalid   (lcl_cl_sh_ddra_q2.rvalid),
    .m_axi_rready   (lcl_cl_sh_ddra_q2.rready)
);

dest_register_slice DDR_A_TST_AXI4_REG_SLC_2 (
    .aclk           (aclk),
    .aresetn        (aresetn),
    .s_axi_awid     (lcl_cl_sh_ddra_q2.awid),
    .s_axi_awaddr   (lcl_cl_sh_ddra_q2.awaddr),
    .s_axi_awlen    (lcl_cl_sh_ddra_q2.awlen),
    .s_axi_awsize   (lcl_cl_sh_ddra_q2.awsize),
    .s_axi_awburst  (2'b1),
    .s_axi_awlock   (1'b0),
    .s_axi_awcache  (4'b11),
    .s_axi_awprot   (3'b10),
    .s_axi_awregion (4'b0),
    .s_axi_awqos    (4'b0),
    .s_axi_awvalid  (lcl_cl_sh_ddra_q2.awvalid),
    .s_axi_awready  (lcl_cl_sh_ddra_q2.awready),
    .s_axi_wdata    (lcl_cl_sh_ddra_q2.wdata),
    .s_axi_wstrb    (lcl_cl_sh_ddra_q2.wstrb),
    .s_axi_wlast    (lcl_cl_sh_ddra_q2.wlast),
    .s_axi_wvalid   (lcl_cl_sh_ddra_q2.wvalid),
    .s_axi_wready   (lcl_cl_sh_ddra_q2.wready),
    .s_axi_bid      (lcl_cl_sh_ddra_q2.bid),
    .s_axi_bresp    (lcl_cl_sh_ddra_q2.bresp),
    .s_axi_bvalid   (lcl_cl_sh_ddra_q2.bvalid),
    .s_axi_bready   (lcl_cl_sh_ddra_q2.bready),
    .s_axi_arid     (lcl_cl_sh_ddra_q2.arid),
    .s_axi_araddr   (lcl_cl_sh_ddra_q2.araddr),
    .s_axi_arlen    (lcl_cl_sh_ddra_q2.arlen),
    .s_axi_arsize   (lcl_cl_sh_ddra_q2.arsize),
    .s_axi_arburst  (2'b1),
    .s_axi_arlock   (1'b0),
    .s_axi_arcache  (4'b11),
    .s_axi_arprot   (3'b10),
    .s_axi_arregion (4'b0),
    .s_axi_arqos    (4'b0),
    .s_axi_arvalid  (lcl_cl_sh_ddra_q2.arvalid),
    .s_axi_arready  (lcl_cl_sh_ddra_q2.arready),
    .s_axi_rid      (lcl_cl_sh_ddra_q2.rid),
    .s_axi_rdata    (lcl_cl_sh_ddra_q2.rdata),
    .s_axi_rresp    (lcl_cl_sh_ddra_q2.rresp),
    .s_axi_rlast    (lcl_cl_sh_ddra_q2.rlast),
    .s_axi_rvalid   (lcl_cl_sh_ddra_q2.rvalid),
    .s_axi_rready   (lcl_cl_sh_ddra_q2.rready),
    
    .m_axi_awid     (lcl_cl_sh_ddra.awid),
    .m_axi_awaddr   (lcl_cl_sh_ddra.awaddr),
    .m_axi_awlen    (lcl_cl_sh_ddra.awlen),
    .m_axi_awsize   (lcl_cl_sh_ddra.awsize),
    .m_axi_awburst  (),
    .m_axi_awlock   (),
    .m_axi_awcache  (),
    .m_axi_awprot   (),
    .m_axi_awregion (),
    .m_axi_awqos    (),
    .m_axi_awvalid  (lcl_cl_sh_ddra.awvalid),
    .m_axi_awready  (lcl_cl_sh_ddra.awready),
    .m_axi_wdata    (lcl_cl_sh_ddra.wdata),
    .m_axi_wstrb    (lcl_cl_sh_ddra.wstrb),
    .m_axi_wlast    (lcl_cl_sh_ddra.wlast),
    .m_axi_wvalid   (lcl_cl_sh_ddra.wvalid),
    .m_axi_wready   (lcl_cl_sh_ddra.wready),
    .m_axi_bid      (lcl_cl_sh_ddra.bid),
    .m_axi_bresp    (lcl_cl_sh_ddra.bresp),
    .m_axi_bvalid   (lcl_cl_sh_ddra.bvalid),
    .m_axi_bready   (lcl_cl_sh_ddra.bready),
    .m_axi_arid     (lcl_cl_sh_ddra.arid),
    .m_axi_araddr   (lcl_cl_sh_ddra.araddr),
    .m_axi_arlen    (lcl_cl_sh_ddra.arlen),
    .m_axi_arsize   (lcl_cl_sh_ddra.arsize),
    .m_axi_arburst  (),
    .m_axi_arlock   (),
    .m_axi_arcache  (),
    .m_axi_arprot   (),
    .m_axi_arregion (),
    .m_axi_arqos    (),
    .m_axi_arvalid  (lcl_cl_sh_ddra.arvalid),
    .m_axi_arready  (lcl_cl_sh_ddra.arready),
    .m_axi_rid      (lcl_cl_sh_ddra.rid),
    .m_axi_rdata    (lcl_cl_sh_ddra.rdata),
    .m_axi_rresp    (lcl_cl_sh_ddra.rresp),
    .m_axi_rlast    (lcl_cl_sh_ddra.rlast),
    .m_axi_rvalid   (lcl_cl_sh_ddra.rvalid),
    .m_axi_rready   (lcl_cl_sh_ddra.rready)
);
//assign lcl_cl_sh_ddra.awid[15:9] = 7'b0;
//assign lcl_cl_sh_ddra.wid[15:9] = 7'b0;
//assign lcl_cl_sh_ddra.arid[15:9] = 7'b0;

//----------------------------
// flop the output of interconnect for DDRB
// back to back for SLR crossing
//----------------------------

//back to back register slices for SLR crossing
src_register_slice DDR_B_TST_AXI4_REG_SLC_1 (
    .aclk           (aclk),
    .aresetn        (aresetn),
    .s_axi_awid     (lcl_cl_sh_ddrb_q.awid),
    .s_axi_awaddr   ({lcl_cl_sh_ddrb_q.awaddr[63:36], 2'b0, lcl_cl_sh_ddrb_q.awaddr[33:0]}),
    .s_axi_awlen    (lcl_cl_sh_ddrb_q.awlen),
    .s_axi_awsize   (lcl_cl_sh_ddrb_q.awsize),
    .s_axi_awburst  (2'b1),
    .s_axi_awlock   (1'b0),
    .s_axi_awcache  (4'b11),
    .s_axi_awprot   (3'b10),
    .s_axi_awregion (4'b0),
    .s_axi_awqos    (4'b0),
    .s_axi_awvalid  (lcl_cl_sh_ddrb_q.awvalid),
    .s_axi_awready  (lcl_cl_sh_ddrb_q.awready),
    .s_axi_wdata    (lcl_cl_sh_ddrb_q.wdata),
    .s_axi_wstrb    (lcl_cl_sh_ddrb_q.wstrb),
    .s_axi_wlast    (lcl_cl_sh_ddrb_q.wlast),
    .s_axi_wvalid   (lcl_cl_sh_ddrb_q.wvalid),
    .s_axi_wready   (lcl_cl_sh_ddrb_q.wready),
    .s_axi_bid      (lcl_cl_sh_ddrb_q.bid),
    .s_axi_bresp    (lcl_cl_sh_ddrb_q.bresp),
    .s_axi_bvalid   (lcl_cl_sh_ddrb_q.bvalid),
    .s_axi_bready   (lcl_cl_sh_ddrb_q.bready),
    .s_axi_arid     (lcl_cl_sh_ddrb_q.arid),
    .s_axi_araddr   ({lcl_cl_sh_ddrb_q.araddr[63:36], 2'b0, lcl_cl_sh_ddrb_q.araddr[33:0]}),
    .s_axi_arlen    (lcl_cl_sh_ddrb_q.arlen),
    .s_axi_arsize   (lcl_cl_sh_ddrb_q.arsize),
    .s_axi_arburst  (2'b1),
    .s_axi_arlock   (1'b0),
    .s_axi_arcache  (4'b11),
    .s_axi_arprot   (3'b10),
    .s_axi_arregion (4'b0),
    .s_axi_arqos    (4'b0),
    .s_axi_arvalid  (lcl_cl_sh_ddrb_q.arvalid),
    .s_axi_arready  (lcl_cl_sh_ddrb_q.arready),
    .s_axi_rid      (lcl_cl_sh_ddrb_q.rid),
    .s_axi_rdata    (lcl_cl_sh_ddrb_q.rdata),
    .s_axi_rresp    (lcl_cl_sh_ddrb_q.rresp),
    .s_axi_rlast    (lcl_cl_sh_ddrb_q.rlast),
    .s_axi_rvalid   (lcl_cl_sh_ddrb_q.rvalid),
    .s_axi_rready   (lcl_cl_sh_ddrb_q.rready),
    
    .m_axi_awid     (lcl_cl_sh_ddrb_q2.awid),
    .m_axi_awaddr   (lcl_cl_sh_ddrb_q2.awaddr),
    .m_axi_awlen    (lcl_cl_sh_ddrb_q2.awlen),
    .m_axi_awsize   (lcl_cl_sh_ddrb_q2.awsize),
    .m_axi_awburst  (),
    .m_axi_awlock   (),
    .m_axi_awcache  (),
    .m_axi_awprot   (),
    .m_axi_awregion (),
    .m_axi_awqos    (),
    .m_axi_awvalid  (lcl_cl_sh_ddrb_q2.awvalid),
    .m_axi_awready  (lcl_cl_sh_ddrb_q2.awready),
    .m_axi_wdata    (lcl_cl_sh_ddrb_q2.wdata),
    .m_axi_wstrb    (lcl_cl_sh_ddrb_q2.wstrb),
    .m_axi_wlast    (lcl_cl_sh_ddrb_q2.wlast),
    .m_axi_wvalid   (lcl_cl_sh_ddrb_q2.wvalid),
    .m_axi_wready   (lcl_cl_sh_ddrb_q2.wready),
    .m_axi_bid      (lcl_cl_sh_ddrb_q2.bid),
    .m_axi_bresp    (lcl_cl_sh_ddrb_q2.bresp),
    .m_axi_bvalid   (lcl_cl_sh_ddrb_q2.bvalid),
    .m_axi_bready   (lcl_cl_sh_ddrb_q2.bready),
    .m_axi_arid     (lcl_cl_sh_ddrb_q2.arid),
    .m_axi_araddr   (lcl_cl_sh_ddrb_q2.araddr),
    .m_axi_arlen    (lcl_cl_sh_ddrb_q2.arlen),
    .m_axi_arsize   (lcl_cl_sh_ddrb_q2.arsize),
    .m_axi_arburst  (),
    .m_axi_arlock   (),
    .m_axi_arcache  (),
    .m_axi_arprot   (),
    .m_axi_arregion (),
    .m_axi_arqos    (),
    .m_axi_arvalid  (lcl_cl_sh_ddrb_q2.arvalid),
    .m_axi_arready  (lcl_cl_sh_ddrb_q2.arready),
    .m_axi_rid      (lcl_cl_sh_ddrb_q2.rid),
    .m_axi_rdata    (lcl_cl_sh_ddrb_q2.rdata),
    .m_axi_rresp    (lcl_cl_sh_ddrb_q2.rresp),
    .m_axi_rlast    (lcl_cl_sh_ddrb_q2.rlast),
    .m_axi_rvalid   (lcl_cl_sh_ddrb_q2.rvalid),
    .m_axi_rready   (lcl_cl_sh_ddrb_q2.rready)
);

dest_register_slice DDR_B_TST_AXI4_REG_SLC_2 (
    .aclk           (aclk),
    .aresetn        (aresetn),
    .s_axi_awid     (lcl_cl_sh_ddrb_q2.awid),
    .s_axi_awaddr   (lcl_cl_sh_ddrb_q2.awaddr),
    .s_axi_awlen    (lcl_cl_sh_ddrb_q2.awlen),
    .s_axi_awsize   (lcl_cl_sh_ddrb_q2.awsize),
    .s_axi_awburst  (2'b1),
    .s_axi_awlock   (1'b0),
    .s_axi_awcache  (4'b11),
    .s_axi_awprot   (3'b10),
    .s_axi_awregion (4'b0),
    .s_axi_awqos    (4'b0),
    .s_axi_awvalid  (lcl_cl_sh_ddrb_q2.awvalid),
    .s_axi_awready  (lcl_cl_sh_ddrb_q2.awready),
    .s_axi_wdata    (lcl_cl_sh_ddrb_q2.wdata),
    .s_axi_wstrb    (lcl_cl_sh_ddrb_q2.wstrb),
    .s_axi_wlast    (lcl_cl_sh_ddrb_q2.wlast),
    .s_axi_wvalid   (lcl_cl_sh_ddrb_q2.wvalid),
    .s_axi_wready   (lcl_cl_sh_ddrb_q2.wready),
    .s_axi_bid      (lcl_cl_sh_ddrb_q2.bid),
    .s_axi_bresp    (lcl_cl_sh_ddrb_q2.bresp),
    .s_axi_bvalid   (lcl_cl_sh_ddrb_q2.bvalid),
    .s_axi_bready   (lcl_cl_sh_ddrb_q2.bready),
    .s_axi_arid     (lcl_cl_sh_ddrb_q2.arid),
    .s_axi_araddr   (lcl_cl_sh_ddrb_q2.araddr),
    .s_axi_arlen    (lcl_cl_sh_ddrb_q2.arlen),
    .s_axi_arsize   (lcl_cl_sh_ddrb_q2.arsize),
    .s_axi_arburst  (2'b1),
    .s_axi_arlock   (1'b0),
    .s_axi_arcache  (4'b11),
    .s_axi_arprot   (3'b10),
    .s_axi_arregion (4'b0),
    .s_axi_arqos    (4'b0),
    .s_axi_arvalid  (lcl_cl_sh_ddrb_q2.arvalid),
    .s_axi_arready  (lcl_cl_sh_ddrb_q2.arready),
    .s_axi_rid      (lcl_cl_sh_ddrb_q2.rid),
    .s_axi_rdata    (lcl_cl_sh_ddrb_q2.rdata),
    .s_axi_rresp    (lcl_cl_sh_ddrb_q2.rresp),
    .s_axi_rlast    (lcl_cl_sh_ddrb_q2.rlast),
    .s_axi_rvalid   (lcl_cl_sh_ddrb_q2.rvalid),
    .s_axi_rready   (lcl_cl_sh_ddrb_q2.rready),
    
    .m_axi_awid     (lcl_cl_sh_ddrb.awid),
    .m_axi_awaddr   (lcl_cl_sh_ddrb.awaddr),
    .m_axi_awlen    (lcl_cl_sh_ddrb.awlen),
    .m_axi_awsize   (lcl_cl_sh_ddrb.awsize),
    .m_axi_awburst  (),
    .m_axi_awlock   (),
    .m_axi_awcache  (),
    .m_axi_awprot   (),
    .m_axi_awregion (),
    .m_axi_awqos    (),
    .m_axi_awvalid  (lcl_cl_sh_ddrb.awvalid),
    .m_axi_awready  (lcl_cl_sh_ddrb.awready),
    .m_axi_wdata    (lcl_cl_sh_ddrb.wdata),
    .m_axi_wstrb    (lcl_cl_sh_ddrb.wstrb),
    .m_axi_wlast    (lcl_cl_sh_ddrb.wlast),
    .m_axi_wvalid   (lcl_cl_sh_ddrb.wvalid),
    .m_axi_wready   (lcl_cl_sh_ddrb.wready),
    .m_axi_bid      (lcl_cl_sh_ddrb.bid),
    .m_axi_bresp    (lcl_cl_sh_ddrb.bresp),
    .m_axi_bvalid   (lcl_cl_sh_ddrb.bvalid),
    .m_axi_bready   (lcl_cl_sh_ddrb.bready),
    .m_axi_arid     (lcl_cl_sh_ddrb.arid),
    .m_axi_araddr   (lcl_cl_sh_ddrb.araddr),
    .m_axi_arlen    (lcl_cl_sh_ddrb.arlen),
    .m_axi_arsize   (lcl_cl_sh_ddrb.arsize),
    .m_axi_arburst  (),
    .m_axi_arlock   (),
    .m_axi_arcache  (),
    .m_axi_arprot   (),
    .m_axi_arregion (),
    .m_axi_arqos    (),
    .m_axi_arvalid  (lcl_cl_sh_ddrb.arvalid),
    .m_axi_arready  (lcl_cl_sh_ddrb.arready),
    .m_axi_rid      (lcl_cl_sh_ddrb.rid),
    .m_axi_rdata    (lcl_cl_sh_ddrb.rdata),
    .m_axi_rresp    (lcl_cl_sh_ddrb.rresp),
    .m_axi_rlast    (lcl_cl_sh_ddrb.rlast),
    .m_axi_rvalid   (lcl_cl_sh_ddrb.rvalid),
    .m_axi_rready   (lcl_cl_sh_ddrb.rready)
);
//assign lcl_cl_sh_ddrb.awid[15:9] = 7'b0;
//assign lcl_cl_sh_ddrb.wid[15:9] = 7'b0;
//assign lcl_cl_sh_ddrb.arid[15:9] = 7'b0;


//----------------------------
// flop the output of interconnect for DDRD
// back to back for SLR crossing
//----------------------------

//back to back register slices for SLR crossing
src_register_slice DDR_D_TST_AXI4_REG_SLC_1 (
    .aclk           (aclk),
    .aresetn        (aresetn),
    .s_axi_awid     (lcl_cl_sh_ddrd_q.awid),
    .s_axi_awaddr   ({lcl_cl_sh_ddrd_q.awaddr[63:36], 2'b0, lcl_cl_sh_ddrd_q.awaddr[33:0]}),
    .s_axi_awlen    (lcl_cl_sh_ddrd_q.awlen),
    .s_axi_awsize   (lcl_cl_sh_ddrd_q.awsize),
    .s_axi_awburst  (2'b1),
    .s_axi_awlock   (1'b0),
    .s_axi_awcache  (4'b11),
    .s_axi_awprot   (3'b10),
    .s_axi_awregion (4'b0),
    .s_axi_awqos    (4'b0),
    .s_axi_awvalid  (lcl_cl_sh_ddrd_q.awvalid),
    .s_axi_awready  (lcl_cl_sh_ddrd_q.awready),
    .s_axi_wdata    (lcl_cl_sh_ddrd_q.wdata),
    .s_axi_wstrb    (lcl_cl_sh_ddrd_q.wstrb),
    .s_axi_wlast    (lcl_cl_sh_ddrd_q.wlast),
    .s_axi_wvalid   (lcl_cl_sh_ddrd_q.wvalid),
    .s_axi_wready   (lcl_cl_sh_ddrd_q.wready),
    .s_axi_bid      (lcl_cl_sh_ddrd_q.bid),
    .s_axi_bresp    (lcl_cl_sh_ddrd_q.bresp),
    .s_axi_bvalid   (lcl_cl_sh_ddrd_q.bvalid),
    .s_axi_bready   (lcl_cl_sh_ddrd_q.bready),
    .s_axi_arid     (lcl_cl_sh_ddrd_q.arid),
    .s_axi_araddr   ({lcl_cl_sh_ddrd_q.araddr[63:36], 2'b0, lcl_cl_sh_ddrd_q.araddr[33:0]}),
    .s_axi_arlen    (lcl_cl_sh_ddrd_q.arlen),
    .s_axi_arsize   (lcl_cl_sh_ddrd_q.arsize),
    .s_axi_arburst  (2'b1),
    .s_axi_arlock   (1'b0),
    .s_axi_arcache  (4'b11),
    .s_axi_arprot   (3'b10),
    .s_axi_arregion (4'b0),
    .s_axi_arqos    (4'b0),
    .s_axi_arvalid  (lcl_cl_sh_ddrd_q.arvalid),
    .s_axi_arready  (lcl_cl_sh_ddrd_q.arready),
    .s_axi_rid      (lcl_cl_sh_ddrd_q.rid),
    .s_axi_rdata    (lcl_cl_sh_ddrd_q.rdata),
    .s_axi_rresp    (lcl_cl_sh_ddrd_q.rresp),
    .s_axi_rlast    (lcl_cl_sh_ddrd_q.rlast),
    .s_axi_rvalid   (lcl_cl_sh_ddrd_q.rvalid),
    .s_axi_rready   (lcl_cl_sh_ddrd_q.rready),
    
    .m_axi_awid     (lcl_cl_sh_ddrd_q2.awid),
    .m_axi_awaddr   (lcl_cl_sh_ddrd_q2.awaddr),
    .m_axi_awlen    (lcl_cl_sh_ddrd_q2.awlen),
    .m_axi_awsize   (lcl_cl_sh_ddrd_q2.awsize),
    .m_axi_awburst  (),
    .m_axi_awlock   (),
    .m_axi_awcache  (),
    .m_axi_awprot   (),
    .m_axi_awregion (),
    .m_axi_awqos    (),
    .m_axi_awvalid  (lcl_cl_sh_ddrd_q2.awvalid),
    .m_axi_awready  (lcl_cl_sh_ddrd_q2.awready),
    .m_axi_wdata    (lcl_cl_sh_ddrd_q2.wdata),
    .m_axi_wstrb    (lcl_cl_sh_ddrd_q2.wstrb),
    .m_axi_wlast    (lcl_cl_sh_ddrd_q2.wlast),
    .m_axi_wvalid   (lcl_cl_sh_ddrd_q2.wvalid),
    .m_axi_wready   (lcl_cl_sh_ddrd_q2.wready),
    .m_axi_bid      (lcl_cl_sh_ddrd_q2.bid),
    .m_axi_bresp    (lcl_cl_sh_ddrd_q2.bresp),
    .m_axi_bvalid   (lcl_cl_sh_ddrd_q2.bvalid),
    .m_axi_bready   (lcl_cl_sh_ddrd_q2.bready),
    .m_axi_arid     (lcl_cl_sh_ddrd_q2.arid),
    .m_axi_araddr   (lcl_cl_sh_ddrd_q2.araddr),
    .m_axi_arlen    (lcl_cl_sh_ddrd_q2.arlen),
    .m_axi_arsize   (lcl_cl_sh_ddrd_q2.arsize),
    .m_axi_arburst  (),
    .m_axi_arlock   (),
    .m_axi_arcache  (),
    .m_axi_arprot   (),
    .m_axi_arregion (),
    .m_axi_arqos    (),
    .m_axi_arvalid  (lcl_cl_sh_ddrd_q2.arvalid),
    .m_axi_arready  (lcl_cl_sh_ddrd_q2.arready),
    .m_axi_rid      (lcl_cl_sh_ddrd_q2.rid),
    .m_axi_rdata    (lcl_cl_sh_ddrd_q2.rdata),
    .m_axi_rresp    (lcl_cl_sh_ddrd_q2.rresp),
    .m_axi_rlast    (lcl_cl_sh_ddrd_q2.rlast),
    .m_axi_rvalid   (lcl_cl_sh_ddrd_q2.rvalid),
    .m_axi_rready   (lcl_cl_sh_ddrd_q2.rready)
);

dest_register_slice DDR_D_TST_AXI4_REG_SLC_2 (
    .aclk           (aclk),
    .aresetn        (aresetn),
    .s_axi_awid     (lcl_cl_sh_ddrd_q2.awid),
    .s_axi_awaddr   (lcl_cl_sh_ddrd_q2.awaddr),
    .s_axi_awlen    (lcl_cl_sh_ddrd_q2.awlen),
    .s_axi_awsize   (lcl_cl_sh_ddrd_q2.awsize),
    .s_axi_awburst  (2'b1),
    .s_axi_awlock   (1'b0),
    .s_axi_awcache  (4'b11),
    .s_axi_awprot   (3'b10),
    .s_axi_awregion (4'b0),
    .s_axi_awqos    (4'b0),
    .s_axi_awvalid  (lcl_cl_sh_ddrd_q2.awvalid),
    .s_axi_awready  (lcl_cl_sh_ddrd_q2.awready),
    .s_axi_wdata    (lcl_cl_sh_ddrd_q2.wdata),
    .s_axi_wstrb    (lcl_cl_sh_ddrd_q2.wstrb),
    .s_axi_wlast    (lcl_cl_sh_ddrd_q2.wlast),
    .s_axi_wvalid   (lcl_cl_sh_ddrd_q2.wvalid),
    .s_axi_wready   (lcl_cl_sh_ddrd_q2.wready),
    .s_axi_bid      (lcl_cl_sh_ddrd_q2.bid),
    .s_axi_bresp    (lcl_cl_sh_ddrd_q2.bresp),
    .s_axi_bvalid   (lcl_cl_sh_ddrd_q2.bvalid),
    .s_axi_bready   (lcl_cl_sh_ddrd_q2.bready),
    .s_axi_arid     (lcl_cl_sh_ddrd_q2.arid),
    .s_axi_araddr   (lcl_cl_sh_ddrd_q2.araddr),
    .s_axi_arlen    (lcl_cl_sh_ddrd_q2.arlen),
    .s_axi_arsize   (lcl_cl_sh_ddrd_q2.arsize),
    .s_axi_arburst  (2'b1),
    .s_axi_arlock   (1'b0),
    .s_axi_arcache  (4'b11),
    .s_axi_arprot   (3'b10),
    .s_axi_arregion (4'b0),
    .s_axi_arqos    (4'b0),
    .s_axi_arvalid  (lcl_cl_sh_ddrd_q2.arvalid),
    .s_axi_arready  (lcl_cl_sh_ddrd_q2.arready),
    .s_axi_rid      (lcl_cl_sh_ddrd_q2.rid),
    .s_axi_rdata    (lcl_cl_sh_ddrd_q2.rdata),
    .s_axi_rresp    (lcl_cl_sh_ddrd_q2.rresp),
    .s_axi_rlast    (lcl_cl_sh_ddrd_q2.rlast),
    .s_axi_rvalid   (lcl_cl_sh_ddrd_q2.rvalid),
    .s_axi_rready   (lcl_cl_sh_ddrd_q2.rready),
    
    .m_axi_awid     (lcl_cl_sh_ddrd.awid),
    .m_axi_awaddr   (lcl_cl_sh_ddrd.awaddr),
    .m_axi_awlen    (lcl_cl_sh_ddrd.awlen),
    .m_axi_awsize   (lcl_cl_sh_ddrd.awsize),
    .m_axi_awburst  (),
    .m_axi_awlock   (),
    .m_axi_awcache  (),
    .m_axi_awprot   (),
    .m_axi_awregion (),
    .m_axi_awqos    (),
    .m_axi_awvalid  (lcl_cl_sh_ddrd.awvalid),
    .m_axi_awready  (lcl_cl_sh_ddrd.awready),
    .m_axi_wdata    (lcl_cl_sh_ddrd.wdata),
    .m_axi_wstrb    (lcl_cl_sh_ddrd.wstrb),
    .m_axi_wlast    (lcl_cl_sh_ddrd.wlast),
    .m_axi_wvalid   (lcl_cl_sh_ddrd.wvalid),
    .m_axi_wready   (lcl_cl_sh_ddrd.wready),
    .m_axi_bid      (lcl_cl_sh_ddrd.bid),
    .m_axi_bresp    (lcl_cl_sh_ddrd.bresp),
    .m_axi_bvalid   (lcl_cl_sh_ddrd.bvalid),
    .m_axi_bready   (lcl_cl_sh_ddrd.bready),
    .m_axi_arid     (lcl_cl_sh_ddrd.arid),
    .m_axi_araddr   (lcl_cl_sh_ddrd.araddr),
    .m_axi_arlen    (lcl_cl_sh_ddrd.arlen),
    .m_axi_arsize   (lcl_cl_sh_ddrd.arsize),
    .m_axi_arburst  (),
    .m_axi_arlock   (),
    .m_axi_arcache  (),
    .m_axi_arprot   (),
    .m_axi_arregion (),
    .m_axi_arqos    (),
    .m_axi_arvalid  (lcl_cl_sh_ddrd.arvalid),
    .m_axi_arready  (lcl_cl_sh_ddrd.arready),
    .m_axi_rid      (lcl_cl_sh_ddrd.rid),
    .m_axi_rdata    (lcl_cl_sh_ddrd.rdata),
    .m_axi_rresp    (lcl_cl_sh_ddrd.rresp),
    .m_axi_rlast    (lcl_cl_sh_ddrd.rlast),
    .m_axi_rvalid   (lcl_cl_sh_ddrd.rvalid),
    .m_axi_rready   (lcl_cl_sh_ddrd.rready)
);

//assign lcl_cl_sh_ddrd.awid[15:9] = 7'b0;
//assign lcl_cl_sh_ddrd.wid[15:9] = 7'b0;
//assign lcl_cl_sh_ddrd.arid[15:9] = 7'b0;

endmodule

